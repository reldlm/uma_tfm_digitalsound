
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Rodrigo Espejo L�pez de los Mozos
-- 
-- Create Date: 12.03.2024 19:08:22
-- Design Name: 
-- Module Name: tfm_ir_coeff_buffer - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- Instance template
--    tfm_ir_coeff_buffer : entity WORK.tfm_ir_coeff_buffer
--        generic map (
--            bits => bits,
--            ir_d_width => ir_d_width,
--            n_rams => n_rams
--        )
--        port map (
--            sysclk => sysclk,
--            reset => reset,
--            start_tick => start_tick,
--            done_tick => ir_done_tick,
--            dout => ir_output
--        );

entity tfm_ir_coeff_buffer is
    Generic (
        bits : INTEGER := 2;
        ir_d_width : INTEGER := 16;
        n_rams : INTEGER := 2
    );
    Port ( 
        sysclk : in STD_LOGIC;
        reset : in STD_LOGIC;
        start_tick : in STD_LOGIC;
        done_tick : out STD_LOGIC;
        dout : out STD_LOGIC_VECTOR ((ir_d_width*n_rams)-1 downto 0)
        );
end tfm_ir_coeff_buffer;

architecture Behavioral of tfm_ir_coeff_buffer is
    -- Memory
    type memory_block is array ((2**bits-1) downto 0) of STD_LOGIC_VECTOR (ir_d_width-1 downto 0);  -- Array type for the memory
    type ir_buffer is array ((n_rams-1) downto 0) of memory_block;
    signal coeff_s : ir_buffer := (
        -- Block 31
        (
            x"0751", x"06cd", x"05ec", x"04ab", 
            x"0360", x"02a7", x"02f4", x"0400", 
            x"051d", x"05b6", x"0597", x"050a", 
            x"0463", x"03ad", x"02d0", x"01ef", 
            x"0160", x"016c", x"01ff", x"02f0", 
            x"0427", x"0566", x"0667", x"0719", 
            x"073c", x"065b", x"047e", x"023c", 
            x"005c", x"ff12", x"fe2f", x"fd93", 
            x"fda4", x"feb0", x"0045", x"0163", 
            x"0160", x"006b", x"ff34", x"fe78", 
            x"fe82", x"ff05", x"ff8f", x"fff9", 
            x"0037", x"0009", x"ff26", x"fddd", 
            x"fd16", x"fd8a", x"ff16", x"00e4", 
            x"0240", x"02d6", x"02cb", x"027c", 
            x"0227", x"01c0", x"0136", x"0089", 
            x"ffb6", x"feea", x"fe76", x"fe79", 
            x"feec", x"ffd1", x"00dc", x"0176", 
            x"012f", x"001e", x"fecd", x"fd6a", 
            x"fc03", x"fb34", x"fb71", x"fc84", 
            x"fe02", x"ff97", x"0112", x"0244", 
            x"0341", x"042b", x"04ad", x"0424", 
            x"028c", x"00aa", x"ff37", x"fe65", 
            x"fe1f", x"fe36", x"fe3c", x"fdd3", 
            x"fd67", x"fdc5", x"feea", x"fff3", 
            x"0031", x"ff8e", x"fe5d", x"fd24", 
            x"fc11", x"fb55", x"fb3b", x"fbd5", 
            x"fcca", x"fd8b", x"fdc3", x"fd94", 
            x"fd48", x"fd01", x"fc94", x"fbfa", 
            x"fb94", x"fbd7", x"fcbe", x"fd8a", 
            x"fd7d", x"fcb7", x"fbef", x"fbab", 
            x"fc04", x"fcc3", x"fdf6", x"ff92", 
            x"011f", x"01e4", x"0155", x"ff9e", 
            x"fdae", x"fc69", x"fbe0", x"fb86", 
            x"faeb", x"fa22", x"f9d7", x"faa1", 
            x"fc70", x"feb0", x"009d", x"01b8", 
            x"01fd", x"0202", x"0289", x"03cd", 
            x"0538", x"05ac", x"04e2", x"03ad", 
            x"02cf", x"0263", x"0213", x"0164", 
            x"0027", x"fe6f", x"fc9a", x"fb41", 
            x"fadc", x"fb49", x"fc04", x"fc92", 
            x"fceb", x"fd52", x"fdc2", x"fded", 
            x"fd83", x"fc79", x"fb12", x"f9c8", 
            x"f91a", x"f926", x"f9bd", x"fa9f", 
            x"fbab", x"fcc5", x"fdcd", x"fe72", 
            x"fe7c", x"fe13", x"fd95", x"fd69", 
            x"fd96", x"fdd7", x"fdd5", x"fd85", 
            x"fd28", x"fcb5", x"fc10", x"fb5a", 
            x"fad0", x"fa93", x"fa9c", x"fade", 
            x"fb60", x"fbe2", x"fbe4", x"fb4e", 
            x"fa84", x"f9ed", x"f9b8", x"f9e2", 
            x"fa8e", x"fbad", x"fcee", x"fe38", 
            x"ff99", x"0119", x"0268", x"0307", 
            x"02c0", x"01d3", x"00c2", x"000b", 
            x"ffe3", x"fff0", x"ffe4", x"ffd0", 
            x"ffd7", x"ffe0", x"ffab", x"ff4d", 
            x"ff53", x"0025", x"0194", x"02ff", 
            x"03f9", x"0476", x"04cd", x"052c", 
            x"0577", x"0574", x"0519", x"04c3", 
            x"04de", x"055f", x"05b8", x"0570", 
            x"04bb", x"0442", x"0439", x"0406", 
            x"032e", x"01dd", x"00b6", x"005b", 
            x"00e3", x"020f", x"0363", x"0452", 
            x"04c6", x"0506", x"057c", x"0640", 
            x"06ef", x"0742", x"076e", x"07bc", 
            x"086b", x"0960", x"0a7d", x"0b94", 
            x"0c07", x"0b28", x"08ef", x"063c", 
            x"0456", x"03dd", x"0462", x"0521", 
            x"058d", x"0583", x"0533", x"04a2", 
            x"03cb", x"02c0", x"01a3", x"00a4", 
            x"ffa7", x"fe67", x"fd0b", x"fc01", 
            x"fb61", x"fb22", x"fb2f", x"fbaa", 
            x"fc9a", x"fdf1", x"ffae", x"01b2", 
            x"039d", x"04ea", x"0553", x"0511", 
            x"04ff", x"05b8", x"0716", x"08b3", 
            x"0a17", x"0b1c", x"0c1a", x"0d40", 
            x"0e0d", x"0dc3", x"0c17", x"09b2", 
            x"07f3", x"079e", x"0820", x"0846", 
            x"0779", x"05fc", x"0441", x"027d", 
            x"00f1", x"0002", x"ffdf", x"0035", 
            x"0097", x"00a2", x"fff8", x"fe9e", 
            x"fd2c", x"fc5a", x"fc38", x"fc36", 
            x"fbc4", x"fb07", x"facc", x"fb8b", 
            x"fd0d", x"fea2", x"ff95", x"ffa2", 
            x"ff34", x"ff1d", x"ffb7", x"0085", 
            x"00dc", x"0075", x"ffa5", x"ff3b", 
            x"ffa2", x"0089", x"0161", x"01cf", 
            x"019e", x"0099", x"fecd", x"fce1", 
            x"fbb6", x"fbbc", x"fca6", x"fd9d", 
            x"fdf0", x"fd40", x"fbd7", x"fa2d", 
            x"f8a4", x"f75f", x"f663", x"f5cd", 
            x"f5e2", x"f6af", x"f7dc", x"f91e", 
            x"fa55", x"fb65", x"fc2e", x"fc3b", 
            x"fb4e", x"fa1a", x"f9a4", x"fa35", 
            x"fb21", x"fbad", x"fbbb", x"fb96", 
            x"fb6b", x"fb49", x"fb50", x"fb86", 
            x"fbdc", x"fc18", x"fc20", x"fc48", 
            x"fcd2", x"fd87", x"fe00", x"fe0a", 
            x"fdaa", x"fd1a", x"fc96", x"fc1e", 
            x"fba3", x"fae6", x"f9ac", x"f84a", 
            x"f7af", x"f866", x"f9f2", x"fb86", 
            x"fcb5", x"fdac", x"fe80", x"fef3", 
            x"fef3", x"fe94", x"fe18", x"fdd9", 
            x"fdf6", x"fe5d", x"ff0d", x"0027", 
            x"01bd", x"0361", x"0463", x"0477", 
            x"0429", x"0421", x"047b", x"04ed", 
            x"0532", x"0560", x"05c6", x"0666", 
            x"06d1", x"06bb", x"0656", x"060b", 
            x"05ee", x"05a3", x"04d8", x"03b3", 
            x"02b9", x"024b", x"0253", x"0282", 
            x"028d", x"0216", x"0114", x"002f", 
            x"0036", x"010a", x"0198", x"011f", 
            x"ffcb", x"fe4d", x"fce8", x"fb62", 
            x"f9e8", x"f8e7", x"f87f", x"f892", 
            x"f8df", x"f947", x"fa0e", x"fb6d", 
            x"fd00", x"fe0b", x"fe06", x"fd4b", 
            x"fcb6", x"fcd5", x"fda3", x"fead", 
            x"ff94", x"0061", x"0120", x"01b9", 
            x"0227", x"028a", x"0319", x"03c0", 
            x"0438", x"044a", x"03ea", x"033e", 
            x"02a8", x"025e", x"01fc", x"00e0", 
            x"ff41", x"fe1d", x"fdf7", x"fe60", 
            x"fe7b", x"fe08", x"fd39", x"fc39", 
            x"fb2f", x"fa56", x"f9ea", x"fa08", 
            x"fa8e", x"fb19", x"fb74", x"fbad", 
            x"fc0b", x"fc93", x"fcd3", x"fca8", 
            x"fc73", x"fc91", x"fcf6", x"fd89", 
            x"fe43", x"ff20", x"0017", x"0110", 
            x"01f3", x"02a4", x"0345", x"0416", 
            x"050f", x"05a7", x"0582", x"04c9", 
            x"03a7", x"01ff", x"ffc4", x"fd5c", 
            x"fb4c", x"f9ca", x"f8ce", x"f847", 
            x"f81d", x"f860", x"f909", x"f9d9", 
            x"fa7b", x"fab7", x"fab0", x"fad0", 
            x"fb6c", x"fc7c", x"fd8c", x"fe62", 
            x"ff67", x"0149", x"0474", x"0857", 
            x"0bc9", x"0def", x"0e9d", x"0e28", 
            x"0d2b", x"0bec", x"0a80", x"0909", 
            x"07c0", x"06e1", x"0676", x"0663", 
            x"0647", x"05a0", x"043b", x"0269", 
            x"00b6", x"ff41", x"fdd7", x"fc8f", 
            x"fba0", x"fb20", x"fb0b", x"fb7b", 
            x"fc8c", x"fe14", x"ff71", x"0022", 
            x"004c", x"002f", x"0011", x"002d", 
            x"00ac", x"0193", x"0256", x"024f", 
            x"01a0", x"0107", x"011a", x"01d0", 
            x"02a6", x"034e", x"03a5", x"03ac", 
            x"03b1", x"03ba", x"033f", x"01d5", 
            x"ffc9", x"fdee", x"fca8", x"fb91", 
            x"fa65", x"f97d", x"f9a9", x"fb62", 
            x"fe1f", x"0077", x"015b", x"00ec", 
            x"fffa", x"ff0f", x"fe1e", x"fcff", 
            x"fc25", x"fc4f", x"fdd4", x"003e", 
            x"02be", x"04b4", x"05f3", x"0696", 
            x"068b", x"058d", x"03a4", x"0150", 
            x"ff57", x"fe44", x"fe2a", x"fe85", 
            x"fea4", x"fe51", x"fda4", x"fcf2", 
            x"fc94", x"fc96", x"fcc7", x"fc9d", 
            x"fb80", x"f98c", x"f7b5", x"f6fc", 
            x"f788", x"f8a6", x"f9c9", x"fb2b", 
            x"fd05", x"fee0", x"002a", x"00f7", 
            x"01c2", x"02b8", x"0390", x"0435", 
            x"04e7", x"05a9", x"0611", x"05ac", 
            x"048e", x"0340", x"022c", x"0173", 
            x"0103", x"00c7", x"00d4", x"0125", 
            x"0181", x"0194", x"0106", x"ffd5", 
            x"fe5b", x"fd1f", x"fc69", x"fc3a", 
            x"fc6c", x"fc9e", x"fcba", x"fd01", 
            x"fdcf", x"ff32", x"00e2", x"0251", 
            x"030e", x"0314", x"028c", x"01fa", 
            x"021b", x"031f", x"0481", x"05a2", 
            x"0638", x"063e", x"05cf", x"04cd", 
            x"0339", x"0198", x"0079", x"fff1", 
            x"ffbc", x"ffaf", x"ffd6", x"003a", 
            x"0045", x"ff46", x"fd8b", x"fc49", 
            x"fc49", x"fd2f", x"fde7", x"fdaa", 
            x"fc88", x"fb72", x"fb38", x"fbae", 
            x"fbe3", x"fb34", x"f9cb", x"f8a8", 
            x"f89d", x"f994", x"faee", x"fbf8", 
            x"fc73", x"fc7f", x"fc54", x"fc26", 
            x"fc5e", x"fd4a", x"feb0", x"ffee", 
            x"00a4", x"00e5", x"00d5", x"006f", 
            x"fff6", x"ffe6", x"0030", x"005f", 
            x"0040", x"ffe0", x"ff87", x"ff8b", 
            x"ffff", x"0091", x"00d2", x"0065", 
            x"ff73", x"feb9", x"fed0", x"ff52", 
            x"ff67", x"fedd", x"fe20", x"fd9a", 
            x"fd51", x"fcfb", x"fca0", x"fcdf", 
            x"fdfb", x"ff53", x"000c", x"ffd2", 
            x"fedb", x"fd90", x"fc7c", x"fc31", 
            x"fccc", x"fda2", x"fe02", x"fde2", 
            x"fde3", x"fe9c", x"fff7", x"0156", 
            x"023e", x"029e", x"02c6", x"031e", 
            x"03af", x"040d", x"03fe", x"03dc", 
            x"03fc", x"0431", x"0438", x"0443", 
            x"04be", x"05bc", x"069f", x"06d5", 
            x"0654", x"056e", x"0490", x"03c8", 
            x"02df", x"01e1", x"014b", x"01a3", 
            x"02b4", x"03a4", x"03af", x"02e6", 
            x"01d3", x"00f9", x"00b3", x"00ef", 
            x"0158", x"01b8", x"0217", x"0244", 
            x"01d7", x"0099", x"feb4", x"fce8", 
            x"fbfd", x"fc3f", x"fd68", x"fef0", 
            x"0064", x"01ae", x"0306", x"048d", 
            x"0608", x"06fb", x"06f3", x"0606", 
            x"04f3", x"047d", x"04e0", x"05ed", 
            x"0708", x"07b7", x"07f6", x"0804", 
            x"082c", x"0868", x"084a", x"07ad", 
            x"06d7", x"0624", x"058a", x"04be", 
            x"03a5", x"0284", x"01b3", x"0163", 
            x"0169", x"0146", x"007c", x"ff02", 
            x"fd63", x"fc19", x"fb19", x"fa5b", 
            x"f9e4", x"f95e", x"f864", x"f75e", 
            x"f716", x"f7eb", x"f96f", x"faa9", 
            x"faef", x"fab1", x"faa5", x"fafb", 
            x"fb7e", x"fbb3", x"fb7e", x"fb5a", 
            x"fb68", x"fb6b", x"fb42", x"fb43", 
            x"fbcc", x"fca7", x"fd63", x"fdff", 
            x"fe8b", x"feef", x"ff02", x"feac", 
            x"fddc", x"fccc", x"fbf8", x"fbbd", 
            x"fbf4", x"fc37", x"fc90", x"fd32", 
            x"fe08", x"fe85", x"fe3e", x"fd80", 
            x"fd1d", x"fdbc", x"ff19", x"005a", 
            x"00e3", x"00c3", x"006f", x"0065", 
            x"00c5", x"0172", x"020c", x"0241", 
            x"022a", x"0213", x"0203", x"01ca", 
            x"017d", x"0158", x"0161", x"016d", 
            x"0172", x"01bd", x"0240", x"02a7", 
            x"02a4", x"023b", x"01dc", x"0251", 
            x"03d4", x"058b", x"0639", x"0548", 
            x"033b", x"0138", x"000a", x"ffc0", 
            x"ffef", x"0032", x"008a", x"013c", 
            x"0245", x"0358", x"041e", x"0446", 
            x"03b0", x"0255", x"0083", x"fefb", 
            x"fe3f", x"fe26", x"fe55", x"fea7", 
            x"ff2f", x"ffde", x"0052", x"005a", 
            x"0051", x"00a2", x"015c", x"0256", 
            x"0361", x"0453", x"04c4", x"0483", 
            x"03b5", x"02d0", x"0259", x"0256", 
            x"0273", x"024a", x"01d3", x"0152", 
            x"016c", x"0284", x"0421", x"0571", 
            x"05f2", x"05bd", x"050e", x"0406", 
            x"02c3", x"01a5", x"00bf", x"ffd6", 
            x"fee5", x"fe32", x"fe29", x"ff05", 
            x"005e", x"015d", x"015d", x"0077", 
            x"ff5f", x"fe99", x"fe32", x"fddf", 
            x"fd49", x"fca4", x"fc84", x"fd4a", 
            x"fec4", x"002b", x"00a7", x"0041", 
            x"ff86", x"fecf", x"fe4a", x"fe18", 
            x"fe8d", x"ffca", x"0186", x"0361", 
            x"04f0", x"05db", x"0619", x"05f9", 
            x"05b5", x"0557", x"04b8", x"03c9", 
            x"02bd", x"01b9", x"0101", x"00c1", 
            x"00a1", x"0016", x"ff1c", x"fe4c", 
            x"fe37", x"fedc", x"ffc2", x"007e", 
            x"00d3", x"00a6", x"0022", x"ffa8", 
            x"ff78", x"ff77", x"ff54", x"ff23"
        ),
        -- Block 30
        (
            x"ff5a", x"0006", x"00ad", x"00b8", 
            x"0018", x"ff61", x"ff25", x"ff4d", 
            x"ff9e", x"0020", x"008e", x"008a", 
            x"fff1", x"ff10", x"fe73", x"fe46", 
            x"fe2f", x"fdda", x"fd58", x"fd07", 
            x"fd0d", x"fd70", x"fe66", x"0035", 
            x"0260", x"03db", x"0428", x"03aa", 
            x"0348", x"0362", x"03a1", x"03a2", 
            x"036e", x"0303", x"0211", x"008b", 
            x"fef4", x"fe63", x"ff58", x"00dc", 
            x"017b", x"00b7", x"ff5a", x"fe2b", 
            x"fd31", x"fc2a", x"fb04", x"f9f3", 
            x"f92f", x"f886", x"f7c2", x"f719", 
            x"f6dd", x"f701", x"f732", x"f735", 
            x"f725", x"f738", x"f79a", x"f87f", 
            x"fa03", x"fc05", x"fe2a", x"ffab", 
            x"000a", x"ffb2", x"ff92", x"0057", 
            x"01b7", x"02dc", x"0337", x"02d3", 
            x"01d9", x"00b2", x"0020", x"009d", 
            x"01df", x"0300", x"0336", x"027e", 
            x"0165", x"0061", x"ff5e", x"fdea", 
            x"fc02", x"fa51", x"f975", x"f94d", 
            x"f918", x"f873", x"f7a1", x"f714", 
            x"f742", x"f84d", x"f9fb", x"fbcf", 
            x"fd56", x"fe59", x"fee3", x"ff14", 
            x"fef7", x"fed7", x"ff0d", x"ff5c", 
            x"ff2e", x"fe46", x"fd18", x"fc32", 
            x"fbd0", x"fb9e", x"fb12", x"fa42", 
            x"f96e", x"f898", x"f7d7", x"f763", 
            x"f756", x"f79c", x"f7df", x"f7f8", 
            x"f841", x"f8d3", x"f94c", x"f97d", 
            x"f9b9", x"fa85", x"fc15", x"fe04", 
            x"ffd8", x"016e", x"02c2", x"0395", 
            x"0392", x"02b1", x"0180", x"00da", 
            x"011b", x"01ed", x"02af", x"0356", 
            x"0448", x"05ac", x"06f7", x"0760", 
            x"06ce", x"05d9", x"0511", x"0479", 
            x"03ba", x"02b7", x"01d2", x"0174", 
            x"0197", x"01cd", x"0193", x"00b9", 
            x"ff67", x"fdf6", x"fc97", x"fb80", 
            x"fb01", x"fb2a", x"fb9c", x"fbf1", 
            x"fc17", x"fc6e", x"fd61", x"fec4", 
            x"0012", x"00db", x"00da", x"004f", 
            x"ffeb", x"002d", x"00d9", x"0128", 
            x"00c6", x"000d", x"ff9f", x"0004", 
            x"0168", x"035d", x"0536", x"0657", 
            x"06be", x"06df", x"06d8", x"0676", 
            x"05d6", x"0554", x"0516", x"04f7", 
            x"0503", x"053e", x"056a", x"0533", 
            x"04a4", x"0418", x"03db", x"0402", 
            x"0492", x"057f", x"065d", x"0694", 
            x"0600", x"04d5", x"0362", x"0208", 
            x"0136", x"00dd", x"00ab", x"00ab", 
            x"00f6", x"0143", x"00e7", x"ff7f", 
            x"fd75", x"fbda", x"fb97", x"fc96", 
            x"fe1b", x"ff73", x"0080", x"0157", 
            x"01c2", x"016e", x"0054", x"ff21", 
            x"fe7f", x"fe58", x"fe49", x"fe69", 
            x"ff10", x"0051", x"01d2", x"0308", 
            x"039c", x"03cb", x"03e6", x"042c", 
            x"04ca", x"05bc", x"0695", x"06fa", 
            x"0702", x"06f6", x"06fd", x"06f9", 
            x"06c0", x"062d", x"0594", x"0512", 
            x"0469", x"0387", x"028d", x"018c", 
            x"00aa", x"ffd2", x"febd", x"fd4c", 
            x"fb75", x"f96a", x"f7aa", x"f6b8", 
            x"f6e4", x"f807", x"f986", x"faf6", 
            x"fc4a", x"fd83", x"fe7c", x"feef", 
            x"ff09", x"ff65", x"0047", x"0178", 
            x"02a4", x"03cc", x"051e", x"06a1", 
            x"080d", x"08d9", x"08a2", x"07a1", 
            x"069b", x"0636", x"06a2", x"0769", 
            x"07ed", x"07e2", x"0734", x"05c4", 
            x"039b", x"0145", x"ff85", x"fec4", 
            x"feec", x"ff70", x"ffb3", x"ff33", 
            x"fdc6", x"fb86", x"f8d2", x"f65b", 
            x"f4c4", x"f433", x"f469", x"f510", 
            x"f5f4", x"f6e1", x"f79d", x"f815", 
            x"f863", x"f893", x"f8b2", x"f946", 
            x"fadb", x"fd32", x"ff77", x"0113", 
            x"020e", x"0282", x"0271", x"023f", 
            x"02ab", x"03b8", x"047c", x"0440", 
            x"032e", x"01f7", x"0133", x"0108", 
            x"012b", x"0109", x"0086", x"001f", 
            x"003b", x"0076", x"fff2", x"fea7", 
            x"fd7d", x"fd20", x"fd65", x"fdc9", 
            x"fe00", x"fe22", x"fe60", x"feb0", 
            x"ff08", x"ff28", x"fec5", x"fdd9", 
            x"fca0", x"fb6b", x"fa6b", x"f9b3", 
            x"f944", x"f90b", x"f8c1", x"f859", 
            x"f82c", x"f846", x"f84e", x"f82f", 
            x"f864", x"f98f", x"fbfb", x"ff4f", 
            x"02c7", x"0591", x"0716", x"0752", 
            x"067f", x"04c1", x"026c", x"002c", 
            x"fe9c", x"fdbd", x"fd59", x"fd32", 
            x"fcf5", x"fc2a", x"fac7", x"f94d", 
            x"f82e", x"f798", x"f79a", x"f81a", 
            x"f8c0", x"f950", x"f9f3", x"faca", 
            x"fb94", x"fbc4", x"fb73", x"fb72", 
            x"fc67", x"fe44", x"0085", x"0283", 
            x"03d6", x"0471", x"046e", x"03ee", 
            x"034c", x"02ca", x"0229", x"0109", 
            x"ffca", x"ff6b", x"0076", x"028a", 
            x"04b7", x"0621", x"063f", x"04e6", 
            x"0270", x"ff81", x"fcc6", x"fb04", 
            x"faab", x"fb6a", x"fc58", x"fcc4", 
            x"fcfa", x"fd71", x"fe15", x"fe95", 
            x"feef", x"ff97", x"0105", x"0312", 
            x"0508", x"0635", x"065f", x"060b", 
            x"060a", x"0698", x"0768", x"07f0", 
            x"083a", x"0908", x"0ac2", x"0ceb", 
            x"0e8f", x"0ee4", x"0df2", x"0c5f", 
            x"0b17", x"0ad4", x"0b8f", x"0c6f", 
            x"0ca6", x"0c0c", x"0ad1", x"0954", 
            x"07f8", x"06e0", x"0617", x"0593", 
            x"0536", x"04df", x"043d", x"0330", 
            x"0203", x"0128", x"00c6", x"00ee", 
            x"01d5", x"0371", x"04fc", x"057b", 
            x"04d6", x"03a6", x"028e", x"01e4", 
            x"0181", x"012b", x"00f3", x"011a", 
            x"01d1", x"02b1", x"02d6", x"01ec", 
            x"009f", x"000a", x"0090", x"0194", 
            x"022c", x"01e2", x"012f", x"00f5", 
            x"015f", x"01c7", x"01a0", x"0102", 
            x"005a", x"fff7", x"ffe8", x"003d", 
            x"00d9", x"019b", x"0259", x"029d", 
            x"01e2", x"0014", x"fdef", x"fc95", 
            x"fcbf", x"fe4f", x"0048", x"0175", 
            x"0190", x"0157", x"016f", x"01b3", 
            x"0193", x"010d", x"00b8", x"010c", 
            x"01e3", x"0283", x"0266", x"01a4", 
            x"007b", x"ff06", x"fd5c", x"fbb6", 
            x"fa84", x"fa30", x"fac7", x"fc2c", 
            x"fddc", x"fec7", x"fe25", x"fc38", 
            x"f9d9", x"f7e1", x"f71c", x"f802", 
            x"fa32", x"fc92", x"fe3b", x"ff2b", 
            x"fff3", x"00d7", x"01a5", x"0228", 
            x"020b", x"0112", x"ff8f", x"fe6b", 
            x"fe3f", x"fe95", x"fe86", x"fd90", 
            x"fc27", x"fb39", x"fb0a", x"fb11", 
            x"fabf", x"fa15", x"f962", x"f8bf", 
            x"f805", x"f73b", x"f6a9", x"f67a", 
            x"f696", x"f6b2", x"f69c", x"f676", 
            x"f692", x"f77a", x"f988", x"fc68", 
            x"ff4c", x"0155", x"020d", x"0206", 
            x"022e", x"02a3", x"02b7", x"0202", 
            x"0129", x"00e1", x"0153", x"0243", 
            x"033b", x"03b7", x"0394", x"02ed", 
            x"020a", x"014e", x"0097", x"ff57", 
            x"fd57", x"fb04", x"f94d", x"f8cd", 
            x"f942", x"f9c1", x"f9d6", x"fa09", 
            x"fadc", x"fbfc", x"fc8c", x"fc34", 
            x"fb97", x"fb6a", x"fb67", x"fad3", 
            x"f997", x"f865", x"f7c1", x"f7a6", 
            x"f7ce", x"f804", x"f855", x"f8d4", 
            x"f93a", x"f977", x"f9fa", x"fb05", 
            x"fc52", x"fd58", x"fdc5", x"fdaa", 
            x"fd7e", x"fda3", x"fe2a", x"fed6", 
            x"ffb7", x"00e1", x"01fd", x"0297", 
            x"02bc", x"02c6", x"02ec", x"033f", 
            x"03ad", x"040f", x"044c", x"0465", 
            x"04a5", x"0570", x"06b6", x"07d0", 
            x"083b", x"07db", x"06d9", x"0595", 
            x"0465", x"039a", x"0364", x"0362", 
            x"02fc", x"01e9", x"0048", x"fe8c", 
            x"fcf5", x"fb70", x"f9ff", x"f8d9", 
            x"f88d", x"f947", x"fa85", x"fbe1", 
            x"fd4e", x"fedf", x"0025", x"0071", 
            x"ffdb", x"ff4d", x"ffb1", x"0119", 
            x"0310", x"0533", x"0739", x"08d3", 
            x"09dd", x"0a3a", x"09d0", x"08db", 
            x"0833", x"088a", x"099a", x"0a58", 
            x"0a40", x"09a5", x"0906", x"0870", 
            x"075f", x"0582", x"032f", x"0117", 
            x"ffa8", x"feca", x"fdff", x"fcef", 
            x"fbd3", x"fb5b", x"fbce", x"fcbf", 
            x"fd6e", x"fd92", x"fd65", x"fd54", 
            x"fd86", x"fdcf", x"fe18", x"fe54", 
            x"fe93", x"ff38", x"0094", x"0253", 
            x"03a8", x"03e7", x"0331", x"026d", 
            x"0262", x"0300", x"03b1", x"03fa", 
            x"03c6", x"0359", x"02d7", x"0226", 
            x"012b", x"0003", x"ff01", x"fe60", 
            x"fe09", x"fd6a", x"fc29", x"fa94", 
            x"f994", x"f9d0", x"faf9", x"fc4c", 
            x"fd59", x"fe71", x"ffed", x"0166", 
            x"020f", x"01df", x"0196", x"01c4", 
            x"0224", x"0231", x"0230", x"02d5", 
            x"0495", x"06d9", x"0870", x"0898", 
            x"0766", x"05a7", x"042b", x"02f7", 
            x"01ab", x"fff1", x"fdcb", x"fbcb", 
            x"fa88", x"fa26", x"fa69", x"fadc", 
            x"fb41", x"fbb7", x"fc41", x"fcb3", 
            x"fce6", x"fcda", x"fccc", x"fcdf", 
            x"fcfb", x"fd32", x"fda1", x"fe00", 
            x"fe47", x"ff00", x"0071", x"01fb", 
            x"02a3", x"0209", x"00e1", x"0036", 
            x"0058", x"00dd", x"0143", x"0132", 
            x"00c5", x"008a", x"00e4", x"01b2", 
            x"026f", x"0273", x"0180", x"fffa", 
            x"fe95", x"fdc6", x"fd7f", x"fdc3", 
            x"feb2", x"0019", x"017c", x"0257", 
            x"0241", x"013d", x"ffc7", x"feac", 
            x"fec1", x"0037", x"0294", x"051f", 
            x"0731", x"0867", x"08d4", x"08a6", 
            x"079d", x"058c", x"02d2", x"0014", 
            x"fdda", x"fc6f", x"fbbc", x"fb87", 
            x"fbca", x"fca0", x"fdb1", x"fe44", 
            x"fe2b", x"fdee", x"fe1e", x"feb7", 
            x"fed7", x"fd8a", x"fafa", x"f85f", 
            x"f6f9", x"f719", x"f805", x"f911", 
            x"fa1d", x"fb5b", x"fcab", x"fde1", 
            x"fefa", x"fffd", x"00ca", x"0170", 
            x"0224", x"030f", x"042f", x"0566", 
            x"0695", x"077e", x"07be", x"0756", 
            x"06bb", x"0668", x"067a", x"066b", 
            x"05a1", x"03fd", x"0220", x"00d4", 
            x"006f", x"00ce", x"0184", x"0218", 
            x"0244", x"0212", x"01ba", x"015a", 
            x"00dc", x"003d", x"ff96", x"ff10", 
            x"feb5", x"fe7a", x"fe76", x"fed9", 
            x"ff96", x"0003", x"ff64", x"fddc", 
            x"fc52", x"fb90", x"fbb8", x"fc87", 
            x"fdb7", x"fef8", x"0018", x"00fc", 
            x"0191", x"019a", x"00d6", x"ff70", 
            x"fdff", x"fd34", x"fd37", x"fdcb", 
            x"fe86", x"ff32", x"ffe7", x"00cd", 
            x"01d1", x"0294", x"02c2", x"025e", 
            x"0201", x"024e", x"0351", x"048e", 
            x"0565", x"0594", x"0586", x"058a", 
            x"05b2", x"05e8", x"05eb", x"056a", 
            x"044a", x"02de", x"0196", x"00ed", 
            x"0109", x"0184", x"01c1", x"01bd", 
            x"01d0", x"0207", x"023d", x"0231", 
            x"01c3", x"00d4", x"ff7a", x"fe24", 
            x"fd4b", x"fd37", x"fdce", x"feb9", 
            x"ff4f", x"ff0a", x"fe07", x"fcc7", 
            x"fb76", x"fa06", x"f8df", x"f8d2", 
            x"fa3d", x"fc71", x"fe9e", x"0066", 
            x"019c", x"0225", x"022c", x"01f7", 
            x"019d", x"0111", x"0061", x"ffd0", 
            x"ff9f", x"fff5", x"00a4", x"013b", 
            x"0145", x"006b", x"fef9", x"fdbf", 
            x"fd6d", x"fde6", x"fe56", x"fdf2", 
            x"fcda", x"fbef", x"fbc0", x"fc25", 
            x"fc97", x"fcc9", x"fcb0", x"fcb8", 
            x"fd76", x"ff2d", x"017a", x"038e", 
            x"0482", x"0419", x"02c2", x"00d6", 
            x"feae", x"fcf6", x"fc71", x"fd33", 
            x"fe8e", x"ffaf", x"0045", x"0099", 
            x"00cf", x"00a7", x"000a", x"ff33", 
            x"fe49", x"fd3d", x"fc3f", x"fbdf", 
            x"fc5a", x"fd4a", x"fdf4", x"fe0c", 
            x"fde2", x"fdbd", x"fdcb", x"fe0b", 
            x"fe58", x"fe68", x"fdf0", x"fcff", 
            x"fbc3", x"fa5d", x"f918", x"f87b"
        ),
        -- Block 29
        (
            x"f905", x"fa99", x"fc54", x"fd28", 
            x"fcd4", x"fbf0", x"fb51", x"fb6d", 
            x"fc08", x"fcab", x"fd11", x"fd20", 
            x"fcf4", x"fce0", x"fd50", x"fe4d", 
            x"ff32", x"ff36", x"fe04", x"fc00", 
            x"fa4a", x"f9e4", x"fadc", x"fc2d", 
            x"fc4e", x"fab7", x"f83f", x"f664", 
            x"f62a", x"f73f", x"f867", x"f887", 
            x"f7ad", x"f6cb", x"f6d0", x"f7b1", 
            x"f8d0", x"f9d0", x"faaa", x"fb32", 
            x"fb28", x"fa58", x"f8fc", x"f7c2", 
            x"f741", x"f788", x"f85a", x"f9b9", 
            x"fb9c", x"fd81", x"fed6", x"ff7c", 
            x"ffea", x"0072", x"00cb", x"006b", 
            x"ff55", x"fdfa", x"fcd3", x"fc19", 
            x"fb78", x"fa91", x"f968", x"f873", 
            x"f842", x"f8dd", x"f9c3", x"fa7d", 
            x"faf3", x"fb75", x"fc6c", x"fdcc", 
            x"ff3c", x"0062", x"00f5", x"011e", 
            x"012d", x"0147", x"0106", x"0027", 
            x"ff30", x"ff1b", x"0051", x"022e", 
            x"0377", x"039c", x"030a", x"026e", 
            x"0206", x"01a1", x"016c", x"0206", 
            x"039e", x"056f", x"0668", x"0624", 
            x"0532", x"044b", x"0388", x"02c1", 
            x"0217", x"01fe", x"02d9", x"044e", 
            x"0563", x"059e", x"0583", x"05d6", 
            x"06a0", x"0775", x"0853", x"0971", 
            x"0ab2", x"0bdd", x"0cbe", x"0d24", 
            x"0d0f", x"0ca4", x"0c39", x"0bfa", 
            x"0bc8", x"0b66", x"0ac1", x"09ec", 
            x"0922", x"0863", x"0797", x"06cc", 
            x"0607", x"0536", x"0435", x"031d", 
            x"025d", x"026a", x"0335", x"0428", 
            x"04d4", x"055f", x"05e5", x"0638", 
            x"0620", x"059a", x"0507", x"04f9", 
            x"05b9", x"072b", x"08ce", x"0a02", 
            x"0a4c", x"09b1", x"08cf", x"082d", 
            x"07ca", x"073a", x"0641", x"0536", 
            x"04c2", x"0554", x"064c", x"069f", 
            x"05f8", x"048d", x"02a0", x"0082", 
            x"fe8e", x"fd3d", x"fd17", x"fe45", 
            x"002c", x"01a6", x"0199", x"ffd7", 
            x"fd44", x"fb22", x"fa48", x"faa1", 
            x"fb72", x"fc04", x"fc31", x"fcb7", 
            x"fe45", x"0050", x"01d4", x"0223", 
            x"0111", x"fedb", x"fc56", x"fab2", 
            x"fa7a", x"fb3a", x"fc36", x"fd2b", 
            x"fe36", x"ff89", x"0130", x"02eb", 
            x"0457", x"04fa", x"0461", x"028d", 
            x"0030", x"feac", x"ff23", x"0142", 
            x"038a", x"0502", x"05af", x"05b9", 
            x"04e2", x"032a", x"0157", x"003f", 
            x"fff4", x"ffe5", x"ff8d", x"fea8", 
            x"fd68", x"fc18", x"faea", x"fa21", 
            x"f9fd", x"fa71", x"fb44", x"fc7d", 
            x"fe67", x"00c4", x"027b", x"02c8", 
            x"01fe", x"0111", x"00d3", x"013f", 
            x"017e", x"00fb", x"002f", x"0038", 
            x"014a", x"0285", x"0339", x"039f", 
            x"0449", x"0597", x"073c", x"0874", 
            x"0881", x"0791", x"06ba", x"068e", 
            x"0663", x"056c", x"03ce", x"023f", 
            x"0131", x"0088", x"ffef", x"fecc", 
            x"fcb5", x"fa3a", x"f849", x"f769", 
            x"f74a", x"f756", x"f776", x"f7fa", 
            x"f8fc", x"fa01", x"fa63", x"fa1c", 
            x"fa0b", x"fad8", x"fc36", x"fd7f", 
            x"fe86", x"ffa4", x"00eb", x"0231", 
            x"031d", x"033f", x"02a7", x"020d", 
            x"0217", x"028f", x"02ac", x"01ec", 
            x"007c", x"fee4", x"fdcd", x"fdb4", 
            x"fe4d", x"fec3", x"fea7", x"fe64", 
            x"fe88", x"fede", x"fed4", x"fe26", 
            x"fcea", x"fb4c", x"f9b7", x"f8ae", 
            x"f8a5", x"f98f", x"fac1", x"fb96", 
            x"fbc2", x"fb54", x"fac6", x"fa8f", 
            x"fae5", x"fba9", x"fc90", x"fd54", 
            x"fdb8", x"fdc6", x"fdd3", x"fe80", 
            x"002f", x"024e", x"03a2", x"033d", 
            x"011b", x"fe11", x"fb59", x"f9b0", 
            x"f8d2", x"f83e", x"f804", x"f898", 
            x"f9da", x"fafa", x"fb62", x"fb1e", 
            x"fa2a", x"f8b7", x"f764", x"f6e3", 
            x"f77c", x"f8e2", x"fa7a", x"fbda", 
            x"fcd9", x"fd29", x"fc89", x"fb41", 
            x"fa4c", x"faa1", x"fc84", x"ff5d", 
            x"01e7", x"033f", x"0391", x"0379", 
            x"035b", x"0359", x"0380", x"03e8", 
            x"0466", x"04c6", x"0557", x"06a0", 
            x"0873", x"0a06", x"0aa3", x"0a25", 
            x"08da", x"070d", x"0523", x"039b", 
            x"028c", x"01b1", x"0131", x"0148", 
            x"01bf", x"0254", x"0306", x"03c2", 
            x"0461", x"04ab", x"0472", x"038e", 
            x"020c", x"0050", x"fedd", x"fdeb", 
            x"fd3e", x"fc9b", x"fc0c", x"fc0c", 
            x"fcc4", x"fdb7", x"fdf8", x"fd05", 
            x"fb57", x"f9e0", x"f940", x"f943", 
            x"f96a", x"f9a6", x"fa55", x"fba5", 
            x"fd5c", x"ff35", x"00cf", x"0206", 
            x"02b1", x"0282", x"0165", x"0000", 
            x"ff41", x"ff54", x"ff8b", x"ff1b", 
            x"fe3e", x"fdee", x"fea5", x"ffee", 
            x"00d0", x"009d", x"ff7f", x"fe6d", 
            x"fe4e", x"ff06", x"ffc9", x"fffc", 
            x"ff74", x"fe66", x"fd06", x"fba6", 
            x"fab6", x"fa23", x"f986", x"f8fa", 
            x"f910", x"f9fb", x"fb45", x"fc6c", 
            x"fd37", x"fdb3", x"fe3d", x"ff35", 
            x"0091", x"0185", x"0160", x"0075", 
            x"ffac", x"ffaa", x"0052", x"0117", 
            x"01a3", x"0203", x"0235", x"01e7", 
            x"0111", x"001b", x"ff78", x"ff34", 
            x"ff06", x"feb2", x"fe91", x"ff09", 
            x"002e", x"019d", x"029b", x"02c4", 
            x"027d", x"0265", x"029b", x"02e7", 
            x"033b", x"03e4", x"0531", x"070c", 
            x"0909", x"0abf", x"0c0b", x"0cea", 
            x"0d42", x"0cfb", x"0c13", x"0ab0", 
            x"090d", x"0739", x"0539", x"0374", 
            x"0249", x"01cb", x"01ec", x"0269", 
            x"0295", x"01fd", x"00d2", x"ff8d", 
            x"fe0f", x"fbfc", x"f9df", x"f8be", 
            x"f90a", x"fa3c", x"fb92", x"fc97", 
            x"fd6e", x"fe89", x"001d", x"01dc", 
            x"0320", x"03b9", x"041f", x"04fa", 
            x"0657", x"07da", x"0945", x"0a65", 
            x"0ad8", x"0a41", x"08ba", x"0703", 
            x"05d0", x"055a", x"053e", x"050a", 
            x"047a", x"035d", x"01b1", x"ff8e", 
            x"fd20", x"fac1", x"f935", x"f90d", 
            x"fa28", x"fbb4", x"fca0", x"fc6e", 
            x"fb5a", x"fa05", x"f916", x"f8d8", 
            x"f960", x"fa80", x"fb9e", x"fc39", 
            x"fc87", x"fd24", x"fe7d", x"003f", 
            x"01b9", x"02a8", x"035a", x"0414", 
            x"0511", x"0627", x"06a6", x"0628", 
            x"0524", x"0454", x"03f7", x"03c8", 
            x"0378", x"031b", x"02e8", x"030f", 
            x"0388", x"03d7", x"0383", x"0288", 
            x"015b", x"0087", x"004c", x"003d", 
            x"ffc5", x"fec6", x"fdaa", x"fd0b", 
            x"fd15", x"fd7c", x"fdfd", x"fe85", 
            x"ff4d", x"0055", x"013a", x"01c7", 
            x"0221", x"02b1", x"03db", x"0577", 
            x"06da", x"075e", x"0678", x"0408", 
            x"00d1", x"fe37", x"fd5f", x"fe3f", 
            x"ff5c", x"ff22", x"fd7e", x"fb7e", 
            x"fa29", x"f9bb", x"f9c6", x"f9b1", 
            x"f9a2", x"fa04", x"fac9", x"fbbd", 
            x"fcab", x"fd77", x"fe03", x"fe16", 
            x"fd62", x"fc10", x"faeb", x"fa9d", 
            x"faf5", x"fb6e", x"fbb7", x"fc0b", 
            x"fcbd", x"fd8d", x"fde7", x"fd64", 
            x"fc50", x"fbac", x"fc70", x"feac", 
            x"0164", x"034a", x"03fd", x"0445", 
            x"04d0", x"0555", x"0515", x"03ee", 
            x"026d", x"0152", x"0114", x"01a6", 
            x"028e", x"030e", x"027d", x"0091", 
            x"fda5", x"fa62", x"f78a", x"f5b7", 
            x"f503", x"f520", x"f5a9", x"f63e", 
            x"f6d1", x"f77e", x"f843", x"f955", 
            x"fae7", x"fcb2", x"fdf1", x"fe23", 
            x"fda9", x"fd39", x"fceb", x"fc5b", 
            x"fb5c", x"fa92", x"fa8b", x"fb38", 
            x"fc4e", x"fd6c", x"fe2a", x"fe28", 
            x"fd2a", x"fb66", x"f967", x"f773", 
            x"f5c2", x"f4a5", x"f469", x"f525", 
            x"f64a", x"f6f1", x"f6c0", x"f618", 
            x"f58e", x"f53a", x"f4fc", x"f4e4", 
            x"f54b", x"f66d", x"f82b", x"fa26", 
            x"fbf3", x"fd11", x"fd19", x"fc10", 
            x"fa9c", x"f9ed", x"fab5", x"fcf1", 
            x"0009", x"02f9", x"04e2", x"0587", 
            x"054c", x"04e5", x"04b7", x"0490", 
            x"03f0", x"02b7", x"0175", x"00fa", 
            x"0130", x"013c", x"009c", x"ff4a", 
            x"fd96", x"fbe1", x"fa9f", x"f9f8", 
            x"f991", x"f8f6", x"f851", x"f83e", 
            x"f8eb", x"f9b2", x"fa11", x"fa82", 
            x"fbe1", x"fe65", x"0123", x"02d4", 
            x"02e5", x"01da", x"00da", x"00bf", 
            x"0157", x"01ab", x"0138", x"0060", 
            x"0030", x"0112", x"01fd", x"01fe", 
            x"0150", x"00e0", x"0150", x"0290", 
            x"0426", x"0567", x"05c6", x"0578", 
            x"0522", x"0507", x"051f", x"059f", 
            x"06e2", x"08ba", x"0a4f", x"0b05", 
            x"0b41", x"0bba", x"0c50", x"0c3d", 
            x"0b19", x"096a", x"0833", x"07f9", 
            x"0862", x"08ba", x"08c2", x"0896", 
            x"0852", x"0842", x"0890", x"08f8", 
            x"0927", x"0916", x"08da", x"084c", 
            x"0709", x"0517", x"031a", x"0155", 
            x"ffaf", x"fe95", x"feba", x"001d", 
            x"01f0", x"0330", x"0363", x"02a9", 
            x"0181", x"00ab", x"006e", x"002e", 
            x"ff41", x"fdba", x"fc56", x"fbb3", 
            x"fbdb", x"fc84", x"fda3", x"ff47", 
            x"0120", x"02ae", x"0392", x"03ec", 
            x"041b", x"03fe", x"0350", x"0249", 
            x"015f", x"00dd", x"00e0", x"0156", 
            x"020a", x"02db", x"040b", x"0600", 
            x"080c", x"087f", x"06dc", x"04d7", 
            x"0438", x"04f2", x"05a8", x"0570", 
            x"04b7", x"0430", x"03e9", x"034e", 
            x"01ff", x"004b", x"fec6", x"fd90", 
            x"fc5e", x"fb51", x"fad2", x"fb53", 
            x"fcfc", x"ffb1", x"02df", x"0594", 
            x"070e", x"073d", x"06a9", x"0619", 
            x"060c", x"0651", x"0611", x"04c0", 
            x"02f8", x"01b8", x"0146", x"0135", 
            x"0138", x"0154", x"01b7", x"0253", 
            x"02c1", x"02cf", x"0285", x"022c", 
            x"01eb", x"016a", x"0021", x"fe0b", 
            x"fbf2", x"facb", x"fafe", x"fc65", 
            x"fe79", x"0095", x"0222", x"02f0", 
            x"0305", x"02ba", x"026d", x"0233", 
            x"0284", x"03ed", x"0631", x"086c", 
            x"09e4", x"0a85", x"0a97", x"0a54", 
            x"09ae", x"0857", x"0645", x"0425", 
            x"0310", x"0351", x"03e3", x"03a9", 
            x"0284", x"00da", x"ff10", x"fd71", 
            x"fc35", x"fb1e", x"f99f", x"f826", 
            x"f79a", x"f7ef", x"f834", x"f7f3", 
            x"f7d3", x"f878", x"f9c4", x"fb37", 
            x"fc61", x"fcf9", x"fd21", x"fd48", 
            x"fda3", x"fdd8", x"fdaa", x"fd96", 
            x"fe1e", x"ff18", x"0013", x"0117", 
            x"0299", x"04af", x"06ad", x"078f", 
            x"0706", x"0598", x"040a", x"02c7", 
            x"01f7", x"0154", x"003c", x"fe76", 
            x"fc96", x"fbc6", x"fc37", x"fca5", 
            x"fc0d", x"fada", x"fa11", x"fa2c", 
            x"fae8", x"fbac", x"fc05", x"fbbb", 
            x"fb0d", x"fa58", x"fa15", x"fa6e", 
            x"fb2d", x"fc0f", x"fd09", x"fddf", 
            x"fdd6", x"fcb4", x"fb80", x"fb7d", 
            x"fc84", x"fd5f", x"fd56", x"fcd5", 
            x"fc6f", x"fc4a", x"fc46", x"fc58", 
            x"fc3c", x"fb9d", x"fabf", x"fa3e", 
            x"fa6b", x"fb41", x"fc6a", x"fd82", 
            x"fe98", x"0003", x"01a9", x"02fd", 
            x"03ae", x"03f2", x"0418", x"03f6", 
            x"033c", x"01e0", x"0048", x"ff0b", 
            x"fe5b", x"fdff", x"fdaf", x"fd5b", 
            x"fd2c", x"fd73", x"fe6a", x"ffaa", 
            x"004f", x"ffaa", x"fdeb", x"fbe0", 
            x"fa11", x"f889", x"f771", x"f740", 
            x"f835", x"fa00", x"fbe6", x"fd51", 
            x"fe2e", x"feb7", x"ff04", x"ff1d", 
            x"ff55", x"000c", x"0132", x"026c", 
            x"036b", x"0408", x"042d", x"03c7", 
            x"0336", x"02ce", x"0222", x"00a5", 
            x"fee5", x"fe11", x"fe6c", x"fefc"
        ),
        -- Block 28
        (
            x"fed3", x"fe13", x"fd77", x"fd68", 
            x"fd89", x"fd31", x"fc08", x"fa87", 
            x"f96b", x"f8df", x"f87c", x"f830", 
            x"f885", x"f9f8", x"fc38", x"fe17", 
            x"fea9", x"fe14", x"fd28", x"fc59", 
            x"fbab", x"fb3c", x"fb7c", x"fcdd", 
            x"ff4a", x"0216", x"0485", x"05f7", 
            x"062a", x"0585", x"04bc", x"0431", 
            x"03de", x"03b0", x"03ca", x"041d", 
            x"049d", x"053a", x"05a1", x"0544", 
            x"03f5", x"0230", x"007c", x"fef3", 
            x"fdaa", x"fd26", x"fdb0", x"fedb", 
            x"ffbf", x"001d", x"00a4", x"01d1", 
            x"0317", x"036b", x"02a6", x"0196", 
            x"0125", x"015b", x"0161", x"00ba", 
            x"0017", x"0059", x"015c", x"0224", 
            x"021c", x"017e", x"00f8", x"0139", 
            x"0254", x"03b4", x"0469", x"03ec", 
            x"02a5", x"0130", x"ffc2", x"fe62", 
            x"fd14", x"fbe5", x"fae9", x"fa4e", 
            x"fa7e", x"fbc8", x"fdc3", x"ff96", 
            x"00c6", x"0180", x"020b", x"0267", 
            x"0240", x"013e", x"ff96", x"fdfd", 
            x"fd38", x"fd92", x"ff19", x"0165", 
            x"03a0", x"04fd", x"057b", x"058a", 
            x"052a", x"042d", x"02c9", x"019c", 
            x"012f", x"0187", x"020a", x"0209", 
            x"016a", x"007a", x"ff92", x"fee7", 
            x"fe42", x"fd6c", x"fcad", x"fc59", 
            x"fc56", x"fc60", x"fc4d", x"fc53", 
            x"fcae", x"fd35", x"fd8a", x"fd8b", 
            x"fd6e", x"fdba", x"fedc", x"00a1", 
            x"01fc", x"01df", x"0023", x"fd8f", 
            x"fb2d", x"f9ab", x"f939", x"f9cd", 
            x"fb61", x"fd77", x"ff32", x"0021", 
            x"008a", x"0102", x"01f0", x"030f", 
            x"03d3", x"043a", x"04bb", x"05b3", 
            x"071c", x"08f1", x"0b1d", x"0d19", 
            x"0e12", x"0d87", x"0bd0", x"09cc", 
            x"083b", x"0763", x"06fe", x"0665", 
            x"0548", x"03fc", x"02d1", x"01b3", 
            x"0062", x"ff06", x"fe2b", x"fde4", 
            x"fdce", x"fdbc", x"fd92", x"fd6d", 
            x"fd57", x"fd60", x"fdb8", x"fe3c", 
            x"feb5", x"ff65", x"00bc", x"02a5", 
            x"044e", x"0515", x"0560", x"05c6", 
            x"0646", x"0663", x"0608", x"05c2", 
            x"05e2", x"0606", x"05cc", x"054b", 
            x"04c2", x"0488", x"04d7", x"0542", 
            x"0512", x"03ed", x"0252", x"013d", 
            x"00e1", x"00df", x"00e0", x"00c9", 
            x"00a8", x"003f", x"ff88", x"fefe", 
            x"feab", x"fe01", x"fcb3", x"fb4e", 
            x"fad0", x"fbc5", x"fde9", x"0053", 
            x"0220", x"02ba", x"0237", x"0142", 
            x"0088", x"0009", x"ff4e", x"fe5f", 
            x"fded", x"fe5a", x"ff36", x"ffc2", 
            x"ff77", x"fe46", x"fc51", x"fa1e", 
            x"f84d", x"f6fb", x"f5f1", x"f53b", 
            x"f528", x"f60c", x"f7cf", x"f9ee", 
            x"fbf5", x"fd71", x"fe19", x"fe1b", 
            x"fdf8", x"fe37", x"fee2", x"ff60", 
            x"fee8", x"fd51", x"fb9c", x"fb16", 
            x"fbf8", x"fd72", x"fec3", x"ffbc", 
            x"007b", x"014e", x"0241", x"02f3", 
            x"02c6", x"0170", x"ff8b", x"fdfb", 
            x"fd1c", x"fcaf", x"fc5c", x"fc03", 
            x"fbd3", x"fbe6", x"fbff", x"fb9e", 
            x"fae0", x"fa74", x"fac9", x"fbb2", 
            x"fc90", x"fcfa", x"fcd1", x"fc0f", 
            x"fb4e", x"fb62", x"fc51", x"fd37", 
            x"fd26", x"fbe7", x"f9f7", x"f83d", 
            x"f7a0", x"f855", x"f991", x"fa4f", 
            x"fa71", x"fa45", x"fa2d", x"fa81", 
            x"fb36", x"fc14", x"fcfb", x"fdc1", 
            x"fe2a", x"fe36", x"fe12", x"fe0c", 
            x"fe2f", x"fe6c", x"feab", x"ff0e", 
            x"ffa2", x"004a", x"00ee", x"017d", 
            x"01e3", x"024b", x"0349", x"0500", 
            x"06d4", x"081e", x"08b4", x"08a2", 
            x"082d", x"07aa", x"0730", x"06c6", 
            x"0663", x"060d", x"05c4", x"053d", 
            x"0421", x"0238", x"ffa8", x"fd47", 
            x"fc25", x"fc5c", x"fcd4", x"fca2", 
            x"fbeb", x"fb5a", x"fb59", x"fc16", 
            x"fd25", x"fe57", x"ffa3", x"006d", 
            x"004d", x"ff88", x"feff", x"ff75", 
            x"00b2", x"021b", x"0394", x"0567", 
            x"0773", x"091a", x"09c1", x"091a", 
            x"0767", x"0511", x"028d", x"0057", 
            x"fefe", x"fec4", x"ff3b", x"ffbe", 
            x"fff8", x"000a", x"0002", x"ff7f", 
            x"fe68", x"fd3b", x"fc8b", x"fc90", 
            x"fd21", x"fe01", x"ff1a", x"0011", 
            x"0070", x"001b", x"ff7b", x"ff11", 
            x"ff2a", x"ffcd", x"00cd", x"022d", 
            x"03e6", x"05c7", x"07af", x"0994", 
            x"0af4", x"0ad4", x"08d2", x"05f4", 
            x"03bb", x"0292", x"019a", x"0039", 
            x"fea3", x"fd84", x"fd68", x"fe2d", 
            x"ff4e", x"0049", x"00a3", x"0035", 
            x"ff0f", x"fd69", x"fbc6", x"fa70", 
            x"f989", x"f950", x"f9dc", x"fb1d", 
            x"fcdc", x"feba", x"007e", x"024b", 
            x"03fc", x"050a", x"04b1", x"02dd", 
            x"00a6", x"ff4a", x"fef5", x"ff08", 
            x"ff07", x"fef6", x"ff0e", x"ff56", 
            x"ff88", x"ff30", x"fe1d", x"fcb6", 
            x"fb76", x"fa82", x"f9f9", x"f9fb", 
            x"fa5a", x"fab2", x"fac8", x"fab9", 
            x"faf2", x"fb98", x"fc3c", x"fc75", 
            x"fc58", x"fc5c", x"fd1e", x"fec7", 
            x"00b7", x"0250", x"0351", x"03f2", 
            x"04a1", x"0577", x"063c", x"068b", 
            x"0653", x"05d2", x"0524", x"048c", 
            x"0498", x"055b", x"0614", x"05e9", 
            x"043f", x"012b", x"fdd4", x"fb94", 
            x"fb12", x"fba9", x"fbf4", x"fb68", 
            x"faeb", x"fb66", x"fcd0", x"fe2f", 
            x"fe1d", x"fc11", x"f8d3", x"f630", 
            x"f5e5", x"f806", x"fb1b", x"fdf4", 
            x"0044", x"0261", x"0445", x"052b", 
            x"047d", x"02dc", x"0190", x"013b", 
            x"0165", x"0141", x"00d4", x"00ea", 
            x"0226", x"0418", x"0564", x"04c3", 
            x"0233", x"ff2a", x"fd75", x"fdaf", 
            x"ff15", x"00ba", x"021f", x"0322", 
            x"03bc", x"038e", x"025f", x"0095", 
            x"ff1a", x"fedc", x"000a", x"01d2", 
            x"038d", x"053f", x"070e", x"08b5", 
            x"0974", x"0907", x"07c4", x"061f", 
            x"0472", x"02ea", x"01de", x"01c0", 
            x"031a", x"05bb", x"087c", x"0a6b", 
            x"0b82", x"0c36", x"0ca0", x"0c79", 
            x"0bb0", x"0a87", x"08e5", x"0691", 
            x"03e8", x"01c1", x"008f", x"000a", 
            x"ffb8", x"ff65", x"fedd", x"fe15", 
            x"fd99", x"fdcb", x"fdf2", x"fcf4", 
            x"fac6", x"f8af", x"f7e9", x"f8bc", 
            x"fa6c", x"fc13", x"fd3f", x"fe0b", 
            x"febe", x"ff20", x"fe9f", x"fd1a", 
            x"fb6c", x"faf2", x"fc4a", x"fed1", 
            x"0192", x"03eb", x"0523", x"0504", 
            x"0423", x"033a", x"02a9", x"0273", 
            x"029e", x"0318", x"035d", x"02ca", 
            x"0155", x"ff87", x"fe21", x"fdba", 
            x"fe0e", x"fe10", x"fcea", x"fad3", 
            x"f8ce", x"f78c", x"f6a6", x"f54f", 
            x"f388", x"f230", x"f1e7", x"f284", 
            x"f36a", x"f441", x"f55a", x"f703", 
            x"f937", x"fb97", x"fd8e", x"fe70", 
            x"fe0d", x"fd51", x"fd64", x"fe7c", 
            x"ffbc", x"0016", x"ff23", x"fd8b", 
            x"fc83", x"fc8e", x"fd14", x"fd2c", 
            x"fca8", x"fc0e", x"fb70", x"fa38", 
            x"f82a", x"f5ee", x"f481", x"f440", 
            x"f49b", x"f48f", x"f393", x"f22a", 
            x"f152", x"f167", x"f1fa", x"f270", 
            x"f2dd", x"f3f1", x"f666", x"fa43", 
            x"fe5f", x"0101", x"0182", x"0127", 
            x"01cd", x"03e8", x"0646", x"07ad", 
            x"0826", x"0892", x"0904", x"08bc", 
            x"073e", x"04dc", x"0259", x"0050", 
            x"ff06", x"fe73", x"fe78", x"fec6", 
            x"ff07", x"ff22", x"ff42", x"ff70", 
            x"ff90", x"ff89", x"ff77", x"ff7f", 
            x"ffaa", x"fff8", x"006a", x"00f2", 
            x"0159", x"0179", x"0162", x"0114", 
            x"0090", x"0022", x"0050", x"015f", 
            x"0301", x"04ba", x"0682", x"08d9", 
            x"0b78", x"0cc3", x"0b59", x"078e", 
            x"0321", x"004f", x"005e", x"02cd", 
            x"05e5", x"0825", x"0928", x"093d", 
            x"084d", x"062d", x"037b", x"013a", 
            x"0024", x"0028", x"010f", x"0296", 
            x"043f", x"0555", x"05a1", x"0585", 
            x"0554", x"0518", x"050b", x"05a9", 
            x"06eb", x"0841", x"0902", x"08aa", 
            x"0758", x"05e7", x"0550", x"05a9", 
            x"0627", x"061c", x"05b1", x"0578", 
            x"056d", x"04e2", x"0386", x"01e3", 
            x"0076", x"ffaf", x"ffe3", x"00af", 
            x"017a", x"0222", x"02d6", x"03a7", 
            x"044f", x"0487", x"046d", x"040d", 
            x"0332", x"0227", x"01e4", x"0325", 
            x"05a9", x"0864", x"0a5e", x"0b54", 
            x"0ba2", x"0b8f", x"0ac5", x"08f2", 
            x"0654", x"0371", x"00d1", x"fee8", 
            x"fe26", x"feac", x"005b", x"02de", 
            x"053f", x"0677", x"0641", x"052d", 
            x"03f7", x"0290", x"0055", x"fd58", 
            x"fadf", x"fa3c", x"fb68", x"fcee", 
            x"fd47", x"fc83", x"fbe8", x"fc0a", 
            x"fbe6", x"fa3d", x"f76f", x"f523", 
            x"f491", x"f543", x"f594", x"f4bd", 
            x"f3b4", x"f417", x"f64d", x"f8e9", 
            x"fa20", x"f9d8", x"f980", x"fa17", 
            x"fb18", x"fb77", x"fb24", x"fae5", 
            x"fb5d", x"fc36", x"fcc0", x"fcd3", 
            x"fcd3", x"fd51", x"fe90", x"0032", 
            x"0167", x"018b", x"010b", x"0112", 
            x"01cc", x"0202", x"00df", x"ff31", 
            x"fe40", x"fe57", x"fedb", x"ff33", 
            x"feec", x"fdd5", x"fc64", x"fb4b", 
            x"fb09", x"fb8f", x"fc6d", x"fd6e", 
            x"fe45", x"feaa", x"fea0", x"fe5b", 
            x"fdcf", x"fca0", x"fae9", x"f98e", 
            x"f956", x"fa82", x"fca1", x"feb4", 
            x"ffd6", x"ffab", x"fe65", x"fcc1", 
            x"fb6f", x"faa2", x"fa48", x"fa2e", 
            x"fa29", x"fa1d", x"fa67", x"fb96", 
            x"fd9a", x"ff96", x"00e1", x"0191", 
            x"01fe", x"023a", x"0229", x"01dd", 
            x"019f", x"0179", x"0116", x"0094", 
            x"006d", x"00be", x"0163", x"025c", 
            x"03a5", x"04c3", x"04ef", x"03ce", 
            x"021e", x"0149", x"025c", x"04eb", 
            x"075c", x"086a", x"082a", x"0769", 
            x"06c3", x"0644", x"058c", x"0458", 
            x"02c0", x"010e", x"ff89", x"fdd6", 
            x"fb93", x"f95e", x"f8b2", x"fa68", 
            x"fd88", x"0040", x"0198", x"0211", 
            x"0306", x"0529", x"07a9", x"0947", 
            x"0977", x"0884", x"0707", x"05f4", 
            x"0611", x"075c", x"08d8", x"09b2", 
            x"09f8", x"09fa", x"09d9", x"094c", 
            x"080f", x"0643", x"0425", x"01fe", 
            x"0018", x"fe85", x"fd27", x"fbef", 
            x"fad7", x"fa07", x"f9bb", x"f9c6", 
            x"f9e1", x"fa20", x"fa96", x"fb47", 
            x"fc76", x"fe41", x"0003", x"00d3", 
            x"0077", x"ffdc", x"ffda", x"0000", 
            x"ffc4", x"ffa1", x"0093", x"02c7", 
            x"054b", x"06ef", x"0776", x"076d", 
            x"078f", x"0835", x"08b7", x"083e", 
            x"069a", x"044c", x"0232", x"011b", 
            x"0135", x"0229", x"035d", x"0431", 
            x"044d", x"0355", x"01ae", x"0083", 
            x"0079", x"00d8", x"00a3", x"ff87", 
            x"fdc9", x"fbe9", x"fa3a", x"f8e7", 
            x"f7e5", x"f6fc", x"f637", x"f5b4", 
            x"f51b", x"f404", x"f2a9", x"f1ea", 
            x"f27f", x"f3f1", x"f529", x"f595", 
            x"f5a0", x"f65a", x"f860", x"fb94", 
            x"ff42", x"023c", x"03ca", x"0491", 
            x"0588", x"067f", x"0690", x"058c", 
            x"046b", x"0432", x"0486", x"047b", 
            x"0412", x"041a", x"0542", x"0748", 
            x"08fc", x"093d", x"07e2", x"05d1", 
            x"03f2", x"0269", x"0157", x"0137", 
            x"01dd", x"0257", x"01f7", x"00ff", 
            x"0029", x"ff9f", x"feca", x"fd35", 
            x"fb21", x"f932", x"f7aa", x"f665", 
            x"f57a", x"f57f", x"f665", x"f722", 
            x"f6f2", x"f630", x"f5ab", x"f5b8", 
            x"f62e", x"f6f6", x"f7f2", x"f8e1"
        ),
        -- Block 27
        (
            x"f9ce", x"fb09", x"fccb", x"feea", 
            x"00d2", x"01f0", x"0207", x"019d", 
            x"017c", x"01ec", x"0250", x"01bc", 
            x"000d", x"fdf7", x"fc3b", x"faee", 
            x"f9d6", x"f8df", x"f81d", x"f77d", 
            x"f725", x"f7a3", x"f91d", x"faaf", 
            x"fb1a", x"fa3e", x"f945", x"f8f8", 
            x"f8ba", x"f7a4", x"f611", x"f552", 
            x"f666", x"f91a", x"fc74", x"ff5a", 
            x"00fc", x"018b", x"01de", x"0247", 
            x"0236", x"0135", x"ff7e", x"fdd0", 
            x"fcec", x"fd5d", x"ff1f", x"0164", 
            x"0333", x"03d0", x"032b", x"0222", 
            x"01b5", x"0257", x"03ad", x"051a", 
            x"0618", x"063c", x"0547", x"039a", 
            x"01f2", x"00d3", x"006b", x"007c", 
            x"00bc", x"00d2", x"009f", x"0060", 
            x"0043", x"000e", x"ff7e", x"fea7", 
            x"fda1", x"fc80", x"fbff", x"fd1b", 
            x"ffa1", x"0250", x"0452", x"05bb", 
            x"06cd", x"074f", x"06bf", x"0500", 
            x"02d5", x"0189", x"022c", x"0482", 
            x"0771", x"0a02", x"0b94", x"0bbd", 
            x"0a92", x"08ce", x"072d", x"05f0", 
            x"04cd", x"03ab", x"02c2", x"01f3", 
            x"00f3", x"0017", x"0013", x"0132", 
            x"02b6", x"0390", x"0323", x"0196", 
            x"ffc9", x"fea8", x"fe7a", x"fee3", 
            x"ff44", x"ff56", x"ff9b", x"00ea", 
            x"0359", x"05f7", x"07e2", x"08da", 
            x"08d2", x"07d5", x"0698", x"0653", 
            x"078e", x"0979", x"0add", x"0b38", 
            x"0ac2", x"0a0b", x"0982", x"095b", 
            x"0950", x"088b", x"0686", x"03a7", 
            x"0102", x"ff92", x"ff50", x"ff3b", 
            x"fe57", x"fcbb", x"fb69", x"fb14", 
            x"fb58", x"fb0f", x"f95b", x"f6b6", 
            x"f478", x"f39b", x"f441", x"f5ef", 
            x"f81f", x"faa9", x"fd76", x"0020", 
            x"0233", x"03c1", x"0568", x"0772", 
            x"0984", x"0b3e", x"0c77", x"0d41", 
            x"0def", x"0ed2", x"0fe2", x"1083", 
            x"1031", x"0f0c", x"0db9", x"0c82", 
            x"0aee", x"08c2", x"0635", x"0366", 
            x"004a", x"fd08", x"f9e4", x"f759", 
            x"f5ed", x"f587", x"f534", x"f402", 
            x"f1e7", x"efb6", x"ee8c", x"eef4", 
            x"f052", x"f170", x"f1b6", x"f1c1", 
            x"f21d", x"f2da", x"f414", x"f631", 
            x"f92e", x"fc68", x"ff2a", x"00d3", 
            x"00f8", x"ffd1", x"fe47", x"fd1d", 
            x"fc85", x"fc50", x"fc56", x"fc7b", 
            x"fcc5", x"fd1e", x"fd77", x"fdac", 
            x"fd74", x"fc7e", x"facc", x"f8ca", 
            x"f749", x"f6d4", x"f6d1", x"f631", 
            x"f4e0", x"f3ed", x"f3db", x"f43c", 
            x"f4e9", x"f651", x"f8a7", x"fb2d", 
            x"fcc7", x"fd1d", x"fcd3", x"fcb8", 
            x"fcea", x"fcfa", x"fc7b", x"fb71", 
            x"fa40", x"f953", x"f903", x"f9af", 
            x"fb91", x"fe35", x"003c", x"006d", 
            x"fea5", x"fc08", x"fa24", x"f96b", 
            x"f939", x"f91e", x"f987", x"fb01", 
            x"fd56", x"ff81", x"005a", x"ffa6", 
            x"fe32", x"fd04", x"fc5e", x"fbf5", 
            x"fbbe", x"fc19", x"fd40", x"feef", 
            x"00c8", x"02b6", x"049f", x"0627", 
            x"0711", x"0756", x"0746", x"0740", 
            x"0706", x"0631", x"0501", x"0436", 
            x"0445", x"04f6", x"05a8", x"05fb", 
            x"05b6", x"04b5", x"0369", x"024c", 
            x"0150", x"fffa", x"fe3a", x"fcc5", 
            x"fc26", x"fc35", x"fc78", x"fccd", 
            x"fd09", x"fcfd", x"fc96", x"fc0c", 
            x"fbb3", x"fbb9", x"fc6d", x"fdc2", 
            x"ff37", x"0049", x"0111", x"021f", 
            x"03be", x"055c", x"05fa", x"054b", 
            x"03f5", x"02df", x"02a7", x"0376", 
            x"0520", x"073a", x"08eb", x"096d", 
            x"08a0", x"0769", x"06bc", x"0675", 
            x"057b", x"0333", x"008e", x"ff40", 
            x"001b", x"0271", x"04fd", x"069e", 
            x"06ea", x"0682", x"0661", x"068b", 
            x"0630", x"04d5", x"02d2", x"0108", 
            x"0003", x"ffaa", x"ffb6", x"0030", 
            x"0146", x"0316", x"0573", x"078d", 
            x"087a", x"07ce", x"05ca", x"0324", 
            x"0111", x"009a", x"01f1", x"0470", 
            x"06f4", x"0858", x"0827", x"0707", 
            x"064e", x"06e9", x"0870", x"0994", 
            x"0999", x"0905", x"0896", x"0856", 
            x"07db", x"06cb", x"0519", x"02e1", 
            x"009b", x"fef3", x"fe94", x"ffd7", 
            x"0237", x"0457", x"0508", x"043b", 
            x"02a9", x"011a", x"ffb8", x"fe8a", 
            x"fdd0", x"fd9f", x"fdd5", x"fe6e", 
            x"ffd1", x"020d", x"047e", x"0612", 
            x"060b", x"0494", x"02d8", x"0248", 
            x"0347", x"0492", x"04c6", x"03f4", 
            x"033b", x"038b", x"04c5", x"05cb", 
            x"057c", x"0364", x"fff0", x"fc6e", 
            x"fa2d", x"f9b1", x"fa9d", x"fc05", 
            x"fd3f", x"fe38", x"feea", x"ff3f", 
            x"ff06", x"fdec", x"fbfb", x"f9a1", 
            x"f776", x"f5d8", x"f4f4", x"f4fa", 
            x"f5ca", x"f714", x"f8fa", x"fb82", 
            x"fde8", x"ff32", x"ff32", x"fec2", 
            x"ff0d", x"002c", x"0152", x"0232", 
            x"0316", x"0433", x"0563", x"0605", 
            x"057c", x"03a8", x"013f", x"ff5e", 
            x"fe97", x"fece", x"ff60", x"ffb0", 
            x"ffa2", x"ff6c", x"ff1f", x"fec1", 
            x"fe5c", x"fda0", x"fc0a", x"f9c8", 
            x"f7f4", x"f7c5", x"f935", x"fb20", 
            x"fc7f", x"fd0b", x"fd33", x"fd40", 
            x"fd2d", x"fd50", x"fe57", x"009e", 
            x"03ac", x"0686", x"0875", x"0917", 
            x"0888", x"0746", x"05ed", x"04a5", 
            x"031b", x"0137", x"ff9c", x"fefa", 
            x"ff33", x"ffba", x"0075", x"01a7", 
            x"032b", x"045d", x"04c0", x"040a", 
            x"0207", x"ff1c", x"fc58", x"faa9", 
            x"fa08", x"fa2e", x"fb85", x"fe9f", 
            x"02d1", x"069b", x"0908", x"0a4b", 
            x"0b01", x"0b49", x"0ac1", x"096b", 
            x"07e4", x"069f", x"057d", x"0423", 
            x"027d", x"00cc", x"ffbc", x"ffc6", 
            x"009a", x"015b", x"0197", x"019d", 
            x"01d1", x"0214", x"01af", x"003e", 
            x"fe6a", x"fd42", x"fd4f", x"fe38", 
            x"ff27", x"ffa2", x"ffc8", x"ffe3", 
            x"ffb2", x"fe5f", x"fbda", x"f957", 
            x"f85f", x"f938", x"facb", x"fc46", 
            x"fd7f", x"fe6c", x"fe81", x"fd3c", 
            x"fac3", x"f801", x"f5cd", x"f43c", 
            x"f308", x"f259", x"f2bb", x"f46b", 
            x"f6a4", x"f811", x"f823", x"f785", 
            x"f6ed", x"f64d", x"f52c", x"f37d", 
            x"f209", x"f16e", x"f1c2", x"f316", 
            x"f563", x"f863", x"fb82", x"fdcf", 
            x"fec4", x"fed4", x"fea9", x"fe70", 
            x"fdf2", x"fcd2", x"fb18", x"f94e", 
            x"f82a", x"f808", x"f8ac", x"f9c6", 
            x"fb1d", x"fc61", x"fd31", x"fd37", 
            x"fc3e", x"fa9a", x"f93d", x"f90e", 
            x"fa40", x"fc32", x"fde8", x"feeb", 
            x"ff5e", x"ff8c", x"ffab", x"ffdb", 
            x"003b", x"00b0", x"007f", x"fedc", 
            x"fc2c", x"fa3e", x"fa71", x"fc56", 
            x"fe52", x"ff6b", x"fff3", x"00a2", 
            x"01ec", x"03be", x"053d", x"05b4", 
            x"056e", x"054f", x"05d7", x"0682", 
            x"0651", x"04c1", x"0260", x"005f", 
            x"ffa7", x"0032", x"0150", x"02aa", 
            x"0455", x"0621", x"0745", x"072b", 
            x"0607", x"04aa", x"03ca", x"0399", 
            x"03df", x"0423", x"0431", x"04ad", 
            x"063f", x"086e", x"0a12", x"0a53", 
            x"0931", x"075a", x"0578", x"03be", 
            x"021e", x"00ee", x"007c", x"006c", 
            x"ffe8", x"fe5f", x"fc1e", x"fa0e", 
            x"f8cb", x"f84f", x"f84b", x"f86d", 
            x"f895", x"f938", x"faca", x"fcfb", 
            x"fe9b", x"feda", x"fe81", x"fecc", 
            x"ff9e", x"ffc0", x"fe71", x"fc8a", 
            x"fbbc", x"fc91", x"fdc8", x"fe71", 
            x"ff2c", x"00a1", x"028f", x"041f", 
            x"04e7", x"0535", x"058d", x"0646", 
            x"0790", x"0912", x"0a59", x"0b1e", 
            x"0b58", x"0b14", x"0a3f", x"0879", 
            x"05dc", x"0333", x"0130", x"0040", 
            x"00a0", x"0203", x"03c6", x"055b", 
            x"062d", x"05fd", x"0507", x"039a", 
            x"0209", x"004d", x"fe5b", x"fcb9", 
            x"fc82", x"fe76", x"01de", x"052b", 
            x"07dc", x"0a9d", x"0d92", x"0fb9", 
            x"1006", x"0e13", x"0aa4", x"076e", 
            x"05d8", x"05ed", x"0658", x"05db", 
            x"04a0", x"03ac", x"0344", x"02e0", 
            x"01f0", x"003f", x"fdeb", x"fbc2", 
            x"fad1", x"fb88", x"fd2f", x"fe9d", 
            x"ff39", x"ff24", x"fec8", x"fe59", 
            x"fdea", x"fdb7", x"fe0b", x"fecb", 
            x"ff67", x"ffea", x"0107", x"02d6", 
            x"048e", x"058a", x"0629", x"0727", 
            x"086b", x"0919", x"08cc", x"0816", 
            x"07c5", x"0803", x"0864", x"088a", 
            x"0862", x"080a", x"07a0", x"06d9", 
            x"055d", x"0356", x"0149", x"ffba", 
            x"fea7", x"fdc0", x"fcd7", x"fc06", 
            x"fb7c", x"fb06", x"fa69", x"f9c1", 
            x"f92f", x"f8ac", x"f877", x"f8f7", 
            x"f9e6", x"fa72", x"fa19", x"f952", 
            x"f902", x"f98c", x"fa9e", x"fb95", 
            x"fbdf", x"fb9e", x"fb84", x"fbbf", 
            x"fb84", x"fa08", x"f7b5", x"f5d2", 
            x"f530", x"f5a0", x"f6a1", x"f7ea", 
            x"f944", x"fa8c", x"fba3", x"fc89", 
            x"fd67", x"fe5c", x"ff42", x"ffad", 
            x"ff35", x"fe04", x"fcf0", x"fc79", 
            x"fc73", x"fc3c", x"fb25", x"f922", 
            x"f6e9", x"f5a4", x"f5f8", x"f78d", 
            x"f932", x"fa28", x"fae0", x"fc1e", 
            x"fdab", x"fed2", x"ff4b", x"ff39", 
            x"feb2", x"fdce", x"fd13", x"fd18", 
            x"fda3", x"fe20", x"fe67", x"feef", 
            x"005a", x"02a0", x"04d1", x"05e0", 
            x"0581", x"0481", x"03e0", x"03be", 
            x"0332", x"0177", x"feed", x"fd10", 
            x"fd24", x"ff10", x"019d", x"034e", 
            x"0329", x"0188", x"ffca", x"fec5", 
            x"fdb0", x"fb5c", x"f82d", x"f625", 
            x"f70d", x"fa82", x"fe5c", x"00b9", 
            x"0153", x"0102", x"0109", x"0252", 
            x"0461", x"05ee", x"0664", x"064f", 
            x"065a", x"068e", x"0664", x"057b", 
            x"0422", x"02b0", x"0115", x"ffbb", 
            x"ff7b", x"009e", x"026a", x"03c9", 
            x"045e", x"0498", x"04e1", x"051c", 
            x"0511", x"04d8", x"0459", x"031f", 
            x"00f5", x"fe87", x"fcf6", x"fce4", 
            x"fdd5", x"fef1", x"ffcc", x"006f", 
            x"0102", x"016c", x"0183", x"0173", 
            x"0173", x"015c", x"00f9", x"007b", 
            x"ffd8", x"fed7", x"fda7", x"fce7", 
            x"fd0b", x"fd7d", x"fd3c", x"fc3e", 
            x"fb85", x"fbda", x"fd06", x"fe0d", 
            x"fdf5", x"fc85", x"fa6b", x"f8f6", 
            x"f946", x"fb55", x"fe12", x"0078", 
            x"022c", x"0313", x"0347", x"0339", 
            x"0377", x"0436", x"051d", x"05eb", 
            x"06c6", x"07a9", x"0832", x"0808", 
            x"073b", x"062e", x"0535", x"040b", 
            x"023a", x"004d", x"ff50", x"ffa6", 
            x"00aa", x"013c", x"00d6", x"ffc0", 
            x"fe5a", x"fc9f", x"fa55", x"f7c2", 
            x"f619", x"f673", x"f88f", x"fb14", 
            x"fcfd", x"fe4d", x"ff4d", x"0014", 
            x"0066", x"0000", x"feb7", x"fcc5", 
            x"fb17", x"fab9", x"fbec", x"fdbc", 
            x"feeb", x"fef0", x"fe4c", x"fdcf", 
            x"fd92", x"fd02", x"fbba", x"fa01", 
            x"f893", x"f810", x"f839", x"f84b", 
            x"f805", x"f7c7", x"f80c", x"f8fb", 
            x"fa1e", x"fb36", x"fc6d", x"fdc8", 
            x"ff03", x"ffb8", x"ffb3", x"fec7", 
            x"fcfe", x"fb03", x"f9f9", x"fa62", 
            x"fbf9", x"fe09", x"ffc7", x"00c9", 
            x"0118", x"00b6", x"fff4", x"ff56", 
            x"ff56", x"0023", x"016a", x"027a", 
            x"02f2", x"02fc", x"030b", x"0337", 
            x"0309", x"0274", x"021a", x"0242", 
            x"0257", x"0197", x"003d", x"ff96", 
            x"006d", x"0233", x"0378", x"0355", 
            x"0250", x"0187", x"012f", x"00ab", 
            x"ff91", x"fe83", x"fe55", x"feac"
        ),
        -- Block 26
        (
            x"fee4", x"feff", x"ff35", x"ff69", 
            x"ff27", x"fe68", x"fe08", x"feb7", 
            x"fff2", x"0109", x"024b", x"0447", 
            x"063f", x"0691", x"04dc", x"0258", 
            x"0033", x"feb2", x"fd89", x"fcdf", 
            x"fd35", x"febf", x"00cf", x"022d", 
            x"01f6", x"004b", x"fe37", x"fc6a", 
            x"faa0", x"f88f", x"f6a3", x"f5e4", 
            x"f6fc", x"f965", x"fc5b", x"ff4b", 
            x"01e2", x"0433", x"061d", x"0752", 
            x"07cf", x"07dc", x"07f9", x"0889", 
            x"094b", x"0989", x"08ee", x"07d9", 
            x"0784", x"08ce", x"0ad6", x"0c07", 
            x"0c16", x"0c1b", x"0cf8", x"0e2c", 
            x"0e81", x"0d92", x"0bc6", x"096f", 
            x"06d3", x"0478", x"02fc", x"0260", 
            x"020a", x"0166", x"006d", x"ff9d", 
            x"ff46", x"ff4f", x"ff1a", x"fe4b", 
            x"fd8b", x"fdd9", x"ff7b", x"0205", 
            x"0499", x"061c", x"05d9", x"048b", 
            x"03e3", x"04cd", x"067c", x"078c", 
            x"0788", x"072f", x"079b", x"08fc", 
            x"0a4f", x"0a62", x"0947", x"0854", 
            x"0845", x"0839", x"06f7", x"04e7", 
            x"03cb", x"0461", x"0593", x"0639", 
            x"0640", x"0612", x"05bd", x"04fa", 
            x"03ac", x"01ff", x"ffef", x"fd92", 
            x"fbac", x"fb25", x"fbdf", x"fcc6", 
            x"fd2f", x"fda5", x"fe8d", x"ff20", 
            x"fe57", x"fc88", x"fb65", x"fbe8", 
            x"fd16", x"fd33", x"fbac", x"f998", 
            x"f86c", x"f848", x"f827", x"f7b7", 
            x"f7d5", x"f937", x"fb0c", x"fc1c", 
            x"fc43", x"fc26", x"fc0f", x"fbaf", 
            x"fb46", x"fb73", x"fc18", x"fc9e", 
            x"fcc9", x"fd12", x"fe1b", x"ffb2", 
            x"0072", x"ff58", x"fcfb", x"fb04", 
            x"fa94", x"fba9", x"fd9c", x"ffb7", 
            x"015f", x"024e", x"02c7", x"035b", 
            x"0402", x"0459", x"0499", x"052d", 
            x"05a5", x"04de", x"027f", x"ff8f", 
            x"fd8d", x"fcf0", x"fd27", x"fda5", 
            x"fe74", x"ff97", x"0001", x"fe64", 
            x"fb06", x"f779", x"f484", x"f17b", 
            x"ee37", x"ec0d", x"ec19", x"edf5", 
            x"f010", x"f137", x"f189", x"f1e2", 
            x"f2d8", x"f40b", x"f4de", x"f5b3", 
            x"f78c", x"fa21", x"fbf1", x"fc86", 
            x"fd25", x"fed9", x"0092", x"0074", 
            x"fe74", x"fca1", x"fcf7", x"ff2c", 
            x"0152", x"0218", x"01fe", x"024b", 
            x"031e", x"032d", x"01a4", x"ff85", 
            x"fec0", x"002c", x"02ae", x"0469", 
            x"045f", x"030b", x"0107", x"fe68", 
            x"fb24", x"f78a", x"f473", x"f2cb", 
            x"f2cd", x"f3d4", x"f4e7", x"f5c5", 
            x"f6e4", x"f86b", x"f9b1", x"fa48", 
            x"fa67", x"fa76", x"fab6", x"fb40", 
            x"fc0d", x"fcce", x"fd2e", x"fd74", 
            x"fe77", x"0037", x"01ab", x"0210", 
            x"0179", x"0055", x"feef", x"fd7e", 
            x"fc15", x"fa9c", x"f8fb", x"f79d", 
            x"f77c", x"f8de", x"fabe", x"fbc5", 
            x"fbd1", x"fc3b", x"fde4", x"ffd7", 
            x"00d1", x"00d9", x"00cc", x"0145", 
            x"0248", x"03a9", x"052c", x"061b", 
            x"05a7", x"0451", x"0395", x"043b", 
            x"05a5", x"06ce", x"0736", x"0684", 
            x"04c6", x"02b6", x"0156", x"0118", 
            x"0171", x"018d", x"0164", x"019b", 
            x"0297", x"03c8", x"040c", x"0305", 
            x"0193", x"009c", x"ffdf", x"fe65", 
            x"fbfd", x"f9a1", x"f85d", x"f817", 
            x"f813", x"f875", x"fa1a", x"fd2c", 
            x"00cf", x"03c3", x"054b", x"057e", 
            x"04b5", x"0380", x"0299", x"027d", 
            x"0372", x"0565", x"0818", x"0b1c", 
            x"0dc3", x"0fa0", x"1102", x"1223", 
            x"1243", x"107a", x"0d29", x"0a30", 
            x"0918", x"0959", x"0940", x"087a", 
            x"0859", x"09be", x"0bca", x"0cf4", 
            x"0cc2", x"0bcb", x"0ad9", x"0a81", 
            x"0ad8", x"0b46", x"0ada", x"0915", 
            x"069c", x"051a", x"05b8", x"07df", 
            x"09f5", x"0ad1", x"0a8a", x"09ed", 
            x"0984", x"0949", x"08de", x"079d", 
            x"051c", x"01e7", x"ff4d", x"fe5f", 
            x"fef6", x"001a", x"0139", x"0291", 
            x"03f6", x"0471", x"0366", x"014e", 
            x"ff3d", x"fdec", x"fd57", x"fd16", 
            x"fd09", x"fd97", x"ff1e", x"01a5", 
            x"046d", x"062e", x"064d", x"0585", 
            x"04d3", x"0482", x"0498", x"0539", 
            x"0653", x"0774", x"0812", x"07f1", 
            x"0765", x"06fd", x"06ce", x"0671", 
            x"0577", x"03f1", x"027b", x"01a8", 
            x"0151", x"00f1", x"0070", x"000e", 
            x"ff87", x"fec4", x"fe7b", x"fee1", 
            x"ff16", x"fe01", x"fb7f", x"f8ae", 
            x"f6ed", x"f6d2", x"f7db", x"f8d1", 
            x"f8cc", x"f808", x"f736", x"f669", 
            x"f5a1", x"f576", x"f6b6", x"f940", 
            x"fbdd", x"fd7c", x"fe49", x"ff22", 
            x"00ae", x"02c0", x"046b", x"04db", 
            x"0457", x"03f7", x"0467", x"050b", 
            x"04cc", x"0371", x"021c", x"01f9", 
            x"02e5", x"03e1", x"0449", x"0421", 
            x"038e", x"0280", x"013c", x"0041", 
            x"ffa1", x"fedb", x"fd88", x"fc2d", 
            x"fbb6", x"fbe2", x"fba8", x"fb26", 
            x"fba1", x"fdbc", x"0025", x"00bc", 
            x"ff0b", x"fca9", x"fb0c", x"fa2a", 
            x"f96d", x"f8d0", x"f898", x"f89f", 
            x"f8af", x"f903", x"fa25", x"fc1c", 
            x"fe1b", x"ff16", x"fea0", x"fd0f", 
            x"faf4", x"f8da", x"f70b", x"f5d2", 
            x"f51d", x"f429", x"f296", x"f158", 
            x"f1a8", x"f3c0", x"f693", x"f8b4", 
            x"f98c", x"f96c", x"f8c0", x"f7c0", 
            x"f6db", x"f66b", x"f66a", x"f698", 
            x"f704", x"f81a", x"f9ba", x"fb14", 
            x"fb8e", x"fb9a", x"fc06", x"fd00", 
            x"fe59", x"ffca", x"011c", x"01e9", 
            x"01e3", x"0166", x"0122", x"011a", 
            x"00cc", x"0000", x"ff09", x"fe31", 
            x"fcfb", x"fb2b", x"f9a1", x"f954", 
            x"fa4e", x"fbd4", x"fd20", x"fdd8", 
            x"fe34", x"fe68", x"fe32", x"fd0c", 
            x"fa83", x"f711", x"f3db", x"f1dd", 
            x"f16c", x"f25c", x"f487", x"f77e", 
            x"fa9c", x"fd26", x"feac", x"ff70", 
            x"0041", x"0197", x"02c6", x"02e1", 
            x"017f", x"ff64", x"fdc8", x"fd60", 
            x"fe29", x"ffb2", x"015e", x"02a1", 
            x"036d", x"040e", x"04bc", x"056b", 
            x"05b3", x"04f2", x"031c", x"0116", 
            x"ffe0", x"fff2", x"0113", x"02ae", 
            x"0446", x"056d", x"05c6", x"057d", 
            x"0517", x"04f7", x"0582", x"06aa", 
            x"0764", x"067f", x"0418", x"0205", 
            x"023f", x"04e5", x"0860", x"0ae4", 
            x"0b63", x"09ce", x"06f4", x"03e3", 
            x"0182", x"004e", x"ffff", x"ffb5", 
            x"fe93", x"fcb6", x"fb5c", x"fb78", 
            x"fc92", x"fd87", x"fd90", x"fcb6", 
            x"fb50", x"f9e0", x"f915", x"f943", 
            x"f9d2", x"f9f2", x"f970", x"f8b9", 
            x"f846", x"f82e", x"f893", x"f9e5", 
            x"fc7c", x"fff7", x"035d", x"05ef", 
            x"0742", x"0756", x"0675", x"0513", 
            x"039c", x"0247", x"0128", x"0093", 
            x"00fd", x"0293", x"04b7", x"05fb", 
            x"0566", x"0350", x"00bb", x"fe86", 
            x"fd32", x"fd0b", x"fdfb", x"ff8a", 
            x"00f2", x"015a", x"0066", x"fec9", 
            x"fdd4", x"fe0e", x"fea4", x"fe6a", 
            x"fdca", x"fe7b", x"00df", x"0343", 
            x"03f2", x"0328", x"0234", x"01c1", 
            x"0117", x"ff55", x"fd14", x"fc2d", 
            x"fdf5", x"01a9", x"04b4", x"04cf", 
            x"0216", x"fed6", x"fceb", x"fbe4", 
            x"fa40", x"f7e1", x"f683", x"f788", 
            x"fa50", x"fd04", x"fe4c", x"fe6b", 
            x"fe8c", x"ff14", x"ff37", x"fe19", 
            x"fc15", x"fb07", x"fc8c", x"0085", 
            x"055a", x"0932", x"0b0c", x"0b3c", 
            x"0adf", x"0abf", x"0ade", x"0aa4", 
            x"0997", x"074f", x"0412", x"012e", 
            x"ffdc", x"ffa1", x"fee0", x"fce9", 
            x"fab0", x"f96a", x"f964", x"fa62", 
            x"fc1a", x"fdf6", x"ff6f", x"0088", 
            x"01a1", x"02b1", x"0334", x"029d", 
            x"009a", x"fdac", x"fb30", x"fa79", 
            x"fb61", x"fcb9", x"fdcf", x"fed7", 
            x"0019", x"012a", x"0182", x"0123", 
            x"0075", x"ffc8", x"ff5f", x"ff75", 
            x"ffec", x"005f", x"000d", x"fe9c", 
            x"fc5e", x"fa09", x"f874", x"f807", 
            x"f853", x"f8b3", x"f8f7", x"f937", 
            x"f9ba", x"fada", x"fcd8", x"ff8b", 
            x"0245", x"0446", x"0581", x"068f", 
            x"07b2", x"089d", x"08c1", x"07d2", 
            x"0624", x"0477", x"03a8", x"043c", 
            x"05fe", x"0872", x"0b0f", x"0cff", 
            x"0d5a", x"0c04", x"09b4", x"0738", 
            x"051a", x"037b", x"01d8", x"ffb9", 
            x"fd85", x"fc48", x"fc7b", x"fd8c", 
            x"fe75", x"fed9", x"ff1a", x"ff6e", 
            x"ffbd", x"0043", x"0127", x"021a", 
            x"02a5", x"02d1", x"0335", x"0462", 
            x"0615", x"06fb", x"0650", x"050c", 
            x"04c6", x"05e7", x"075b", x"0821", 
            x"0862", x"08b1", x"0902", x"08f0", 
            x"083f", x"0701", x"0573", x"038b", 
            x"015f", x"ff4c", x"fdfd", x"fe49", 
            x"004b", x"02fe", x"04b3", x"0446", 
            x"0252", x"00d5", x"0110", x"024d", 
            x"02b4", x"0189", x"0037", x"00ae", 
            x"0333", x"065f", x"08c1", x"0a3b", 
            x"0b7d", x"0c98", x"0d01", x"0c6b", 
            x"0b40", x"0a3b", x"09dc", x"0a35", 
            x"0b5d", x"0cf3", x"0dcd", x"0ce2", 
            x"0a5b", x"0760", x"0532", x"041e", 
            x"034a", x"01d0", x"ffff", x"ff60", 
            x"00fa", x"03c7", x"05d2", x"0644", 
            x"05eb", x"05be", x"058e", x"04d6", 
            x"03f1", x"0411", x"05a2", x"0797", 
            x"08d0", x"090d", x"089e", x"07fb", 
            x"0795", x"07a6", x"07de", x"07b8", 
            x"0763", x"0796", x"0846", x"0833", 
            x"0680", x"03b0", x"0112", x"ff61", 
            x"fe76", x"fdba", x"fcba", x"fc0b", 
            x"fcd5", x"fef6", x"0096", x"0053", 
            x"fecd", x"fd69", x"fc88", x"fba9", 
            x"fad5", x"fa7a", x"fa9c", x"fb30", 
            x"fc43", x"fd52", x"fd23", x"fb27", 
            x"f877", x"f71c", x"f82c", x"fa7c", 
            x"fba2", x"fa77", x"f851", x"f75d", 
            x"f81a", x"f943", x"f9dd", x"fa46", 
            x"fb19", x"fbdc", x"fb95", x"f9ad", 
            x"f686", x"f32a", x"f0a5", x"efa9", 
            x"efc1", x"efed", x"f007", x"f0c1", 
            x"f278", x"f48b", x"f5b7", x"f54e", 
            x"f3ef", x"f2ad", x"f204", x"f1d9", 
            x"f1c0", x"f165", x"f0c2", x"f017", 
            x"f024", x"f1c4", x"f4a7", x"f710", 
            x"f79c", x"f669", x"f4ca", x"f3e8", 
            x"f3ea", x"f494", x"f5c6", x"f73e", 
            x"f8ba", x"fa01", x"faa3", x"fa17", 
            x"f88a", x"f6e3", x"f5f5", x"f5d0", 
            x"f61f", x"f6cc", x"f79d", x"f843", 
            x"f8c9", x"f98f", x"faf1", x"fcd5", 
            x"fe46", x"fe07", x"fbe6", x"f8ca", 
            x"f5c6", x"f342", x"f112", x"ef4c", 
            x"ee76", x"ef1a", x"f13d", x"f452", 
            x"f76b", x"f9e3", x"fb77", x"fc01", 
            x"fb60", x"f9dd", x"f88e", x"f8a3", 
            x"fa2e", x"fc10", x"fd76", x"fe55", 
            x"ff20", x"ffe9", x"0040", x"fffa", 
            x"ff71", x"ffa5", x"0142", x"03a7", 
            x"057d", x"05e7", x"04da", x"0305", 
            x"0114", x"ff5c", x"fe50", x"fe98", 
            x"0062", x"02b5", x"03f9", x"03cc", 
            x"037b", x"046d", x"06cb", x"0969", 
            x"0a7e", x"08d4", x"04f4", x"00f7", 
            x"fefe", x"ff4a", x"0058", x"00c7", 
            x"00c6", x"00f8", x"0167", x"022b", 
            x"03b4", x"05dd", x"07c8", x"08ed", 
            x"098c", x"0a0b", x"0a31", x"09ca", 
            x"0923", x"0881", x"07b8", x"0669", 
            x"04b9", x"0394", x"0450", x"0742", 
            x"0ada", x"0ccb", x"0c28", x"09fb", 
            x"07c3", x"0624", x"04e7", x"0419", 
            x"044e", x"059f", x"072b", x"0810", 
            x"0841", x"0811", x"078c", x"069a", 
            x"055e", x"0476", x"0466", x"04e2"
        ),
        -- Block 25
        (
            x"0500", x"0432", x"02c4", x"0185", 
            x"00dd", x"0044", x"feec", x"fd43", 
            x"fd0b", x"ff25", x"0218", x"03c1", 
            x"03fe", x"0470", x"05f0", x"0773", 
            x"07b1", x"06b8", x"0581", x"04e7", 
            x"0500", x"0585", x"0629", x"066b", 
            x"05f3", x"052e", x"04c8", x"04f7", 
            x"0590", x"060d", x"05cb", x"0485", 
            x"02d0", x"0166", x"003f", x"fede", 
            x"fd08", x"faf9", x"f93d", x"f845", 
            x"f858", x"f9a2", x"fbb2", x"fdb6", 
            x"fedf", x"fec7", x"fddd", x"fd6b", 
            x"fe86", x"00d2", x"02c9", x"0365", 
            x"02e6", x"022c", x"020d", x"02f0", 
            x"047d", x"05e4", x"06d8", x"07a2", 
            x"088b", x"090c", x"0891", x"0745", 
            x"05f5", x"0534", x"04f8", x"04c8", 
            x"0474", x"0486", x"0543", x"05f3", 
            x"05b5", x"0442", x"0209", x"ffcb", 
            x"fe1b", x"fd4b", x"fd3a", x"fd3d", 
            x"fcf4", x"fc9d", x"fcca", x"fd92", 
            x"fe30", x"fdc4", x"fc1d", x"f9e7", 
            x"f8ab", x"f949", x"fabc", x"fba2", 
            x"fbe7", x"fc75", x"fddc", x"ff97", 
            x"00c0", x"0160", x"0207", x"02cb", 
            x"032d", x"02f3", x"0299", x"02bf", 
            x"036a", x"040f", x"040c", x"0312", 
            x"014d", x"ff25", x"fd48", x"fcab", 
            x"fddc", x"0013", x"01b2", x"0204", 
            x"0193", x"0115", x"00c3", x"008c", 
            x"006b", x"0056", x"003a", x"004c", 
            x"00e8", x"01af", x"01de", x"0190", 
            x"018e", x"01fd", x"0202", x"00e6", 
            x"feb7", x"fbf8", x"f9f9", x"fa21", 
            x"fc27", x"fe25", x"fe64", x"fd04", 
            x"fb79", x"fa7b", x"f9d6", x"f94f", 
            x"f8f1", x"f8bc", x"f8c7", x"f944", 
            x"fa0b", x"fa95", x"fa93", x"fa31", 
            x"f9aa", x"f931", x"f916", x"f94c", 
            x"f90e", x"f7ae", x"f571", x"f347", 
            x"f1ef", x"f16e", x"f1dc", x"f3b3", 
            x"f654", x"f804", x"f799", x"f5d8", 
            x"f4e5", x"f60a", x"f841", x"f996", 
            x"f93c", x"f7f3", x"f6af", x"f5d5", 
            x"f5b3", x"f685", x"f7f3", x"f8d5", 
            x"f872", x"f7a1", x"f7e6", x"f97a", 
            x"fb4d", x"fc8e", x"fd46", x"fdb7", 
            x"fe2c", x"fee8", x"fff9", x"010c", 
            x"01d2", x"0231", x"0214", x"0153", 
            x"0028", x"ff2f", x"fece", x"fef5", 
            x"ff51", x"ff9b", x"ffd9", x"00c8", 
            x"0317", x"0602", x"07ca", x"07b9", 
            x"0699", x"0541", x"039e", x"0154", 
            x"ff04", x"fddf", x"fe43", x"ffad", 
            x"01cb", x"0496", x"0787", x"0986", 
            x"0989", x"0758", x"0447", x"01dc", 
            x"009d", x"005f", x"011e", x"02db", 
            x"050d", x"06fb", x"0802", x"07c7", 
            x"06bb", x"05ca", x"0544", x"04cc", 
            x"0466", x"04d5", x"06c0", x"09af", 
            x"0c4c", x"0dba", x"0e1c", x"0e02", 
            x"0de7", x"0e11", x"0e5f", x"0e64", 
            x"0dfb", x"0d8d", x"0dba", x"0e84", 
            x"0f53", x"0f84", x"0eb3", x"0cf5", 
            x"0b0f", x"09ed", x"098e", x"08d9", 
            x"072e", x"0577", x"0517", x"060f", 
            x"0716", x"06ed", x"051f", x"026e", 
            x"0085", x"007a", x"0171", x"0175", 
            x"ffb2", x"fd8e", x"fd23", x"ff6f", 
            x"03a0", x"07d5", x"0a80", x"0afb", 
            x"09d1", x"0836", x"06c9", x"0593", 
            x"04c4", x"0460", x"0459", x"0493", 
            x"04c9", x"04a4", x"041d", x"035f", 
            x"02ce", x"0242", x"00fc", x"feae", 
            x"fc64", x"fbcc", x"fd63", x"ffc7", 
            x"00e2", x"ffe3", x"fd4a", x"f9e4", 
            x"f649", x"f35a", x"f21a", x"f279", 
            x"f388", x"f4d5", x"f660", x"f7f4", 
            x"f964", x"fae2", x"fc82", x"fdb5", 
            x"fdf6", x"fdcc", x"fe4b", x"ffbf", 
            x"013d", x"0209", x"028b", x"03c2", 
            x"060c", x"08bf", x"0a7c", x"0a25", 
            x"0815", x"05d6", x"042a", x"026e", 
            x"ffce", x"fc6d", x"f944", x"f728", 
            x"f61e", x"f583", x"f484", x"f2e6", 
            x"f161", x"f0b9", x"f111", x"f1de", 
            x"f285", x"f2e3", x"f338", x"f327", 
            x"f1eb", x"efa3", x"eda3", x"ed77", 
            x"ef83", x"f292", x"f513", x"f67b", 
            x"f75e", x"f867", x"f9bc", x"fb53", 
            x"fcd7", x"fe0d", x"ff5d", x"0179", 
            x"044c", x"06ff", x"08cf", x"09b6", 
            x"0a05", x"0986", x"07d2", x"0533", 
            x"0303", x"026c", x"02cf", x"028c", 
            x"0124", x"ffdc", x"0007", x"0163", 
            x"028b", x"02f3", x"0327", x"03db", 
            x"0539", x"0633", x"0551", x"0278", 
            x"ff33", x"fd57", x"fd8a", x"feba", 
            x"ff67", x"fed4", x"fd10", x"fb0d", 
            x"fa15", x"facf", x"fcfa", x"ff6b", 
            x"00c2", x"00c5", x"0028", x"ff7a", 
            x"fead", x"fdb4", x"fd19", x"fd39", 
            x"fdbe", x"fe4a", x"fe91", x"fe79", 
            x"fe83", x"ff89", x"01b0", x"03c9", 
            x"0454", x"0365", x"02b5", x"0370", 
            x"04fe", x"05e9", x"0585", x"04b2", 
            x"04bb", x"05be", x"06db", x"07b6", 
            x"08ba", x"09e3", x"0a32", x"093c", 
            x"07fc", x"07af", x"0860", x"090f", 
            x"08f1", x"07dc", x"05a9", x"0245", 
            x"fea5", x"fc11", x"fae9", x"fa41", 
            x"f934", x"f80d", x"f7d4", x"f8fc", 
            x"fafb", x"fcfd", x"fe75", x"ff36", 
            x"ff54", x"feda", x"fdc0", x"fc09", 
            x"fa0d", x"f8dd", x"f9e6", x"fd63", 
            x"01a7", x"04bd", x"0667", x"07b6", 
            x"093e", x"0a41", x"09a0", x"073e", 
            x"0429", x"018b", x"0010", x"0000", 
            x"0129", x"0302", x"047a", x"0491", 
            x"0375", x"0242", x"0184", x"00dc", 
            x"ff6c", x"fc80", x"f88e", x"f531", 
            x"f3e9", x"f510", x"f7e2", x"fb35", 
            x"fe5e", x"00f7", x"022d", x"0193", 
            x"000e", x"ff16", x"ff45", x"0050", 
            x"0203", x"040e", x"05d5", x"06b7", 
            x"0682", x"0581", x"0422", x"0266", 
            x"0036", x"fdf8", x"fc49", x"fb7f", 
            x"fbc6", x"fce6", x"fdd5", x"fd6b", 
            x"fb64", x"f845", x"f485", x"f035", 
            x"ebd0", x"e8b0", x"e81f", x"ea63", 
            x"eebd", x"f3f9", x"f8cc", x"fc0b", 
            x"fda0", x"fecc", x"00a7", x"02db", 
            x"042d", x"040f", x"0359", x"0381", 
            x"04ed", x"067b", x"069f", x"04be", 
            x"01d9", x"ffa1", x"ff3d", x"0066", 
            x"0191", x"0152", x"ff8a", x"fd0c", 
            x"fabb", x"f8e1", x"f795", x"f72e", 
            x"f7c0", x"f890", x"f8d7", x"f8df", 
            x"f97a", x"facc", x"fb9b", x"fa9b", 
            x"f83d", x"f6d5", x"f836", x"fb9a", 
            x"fef1", x"011d", x"023d", x"02ad", 
            x"0255", x"0107", x"ff2b", x"fd9e", 
            x"fd04", x"fd10", x"fcb8", x"fb64", 
            x"f991", x"f862", x"f8d2", x"faad", 
            x"fc8a", x"fcdb", x"fb58", x"f980", 
            x"f8f5", x"f9d6", x"faea", x"fb2b", 
            x"faca", x"fa63", x"fa02", x"f92e", 
            x"f7f9", x"f751", x"f7e6", x"f93d", 
            x"fa96", x"fc72", x"fff4", x"0487", 
            x"0789", x"06fd", x"0406", x"016d", 
            x"00b3", x"0172", x"0256", x"02a0", 
            x"02f1", x"0466", x"070e", x"099c", 
            x"0aa5", x"09ff", x"08b0", x"0780", 
            x"06e3", x"070e", x"073d", x"0699", 
            x"051c", x"039b", x"02ff", x"0306", 
            x"02e3", x"027a", x"023a", x"0292", 
            x"0387", x"048e", x"04e2", x"0392", 
            x"00b0", x"fdea", x"fd19", x"fe86", 
            x"0116", x"0354", x"042c", x"038a", 
            x"0218", x"00b9", x"ffef", x"ffa1", 
            x"ff36", x"fe09", x"fc2b", x"fa5d", 
            x"f91d", x"f82d", x"f790", x"f7e0", 
            x"f981", x"fbbb", x"fd32", x"fd7b", 
            x"fd89", x"fed5", x"0218", x"065f", 
            x"099d", x"0aaf", x"0ab4", x"0b8d", 
            x"0d58", x"0eb7", x"0f00", x"0ec7", 
            x"0e7f", x"0dd7", x"0c27", x"090e", 
            x"04a9", x"ffa4", x"fb54", x"f91a", 
            x"f91e", x"fa3c", x"fb82", x"fcdf", 
            x"fe5d", x"ff4a", x"fec2", x"fcf8", 
            x"fb1c", x"fa06", x"f92b", x"f792", 
            x"f583", x"f47a", x"f5ba", x"f8f2", 
            x"fc40", x"fda4", x"fccf", x"fb93", 
            x"fbf1", x"fdeb", x"ff8f", x"ffae", 
            x"ff6c", x"00a9", x"0383", x"0637", 
            x"06fb", x"055c", x"027c", x"0011", 
            x"ff2a", x"ff37", x"ff16", x"fee3", 
            x"ffbd", x"01e7", x"03f9", x"04a3", 
            x"047a", x"0485", x"047e", x"03bf", 
            x"0296", x"01eb", x"0256", x"03c7", 
            x"05c9", x"0756", x"0759", x"05f4", 
            x"04a9", x"04e7", x"0707", x"0a38", 
            x"0d2e", x"0f2f", x"108a", x"11b4", 
            x"12a0", x"1314", x"1343", x"1330", 
            x"121b", x"0eed", x"09a6", x"0469", 
            x"01ae", x"01fa", x"03cc", x"0553", 
            x"0630", x"06e7", x"072b", x"05e1", 
            x"0314", x"0093", x"ffc6", x"0005", 
            x"0038", x"0079", x"01a3", x"03e6", 
            x"0665", x"084b", x"0953", x"0946", 
            x"0812", x"0621", x"0401", x"01dc", 
            x"ffc5", x"fe6e", x"fe77", x"ff7c", 
            x"0049", x"ffeb", x"feb0", x"fdc7", 
            x"fdbb", x"fe25", x"fe6b", x"fe00", 
            x"fca6", x"fb37", x"fb58", x"fdba", 
            x"0118", x"0346", x"0354", x"021d", 
            x"0127", x"0135", x"01bb", x"01ac", 
            x"009d", x"ff30", x"fe94", x"ff45", 
            x"0053", x"00a3", x"fff3", x"ff23", 
            x"ff55", x"0088", x"01b9", x"0222", 
            x"0200", x"01b7", x"0122", x"ffd2", 
            x"fe3e", x"fd9a", x"fe2e", x"ff6c", 
            x"0118", x"034d", x"05c6", x"0818", 
            x"09d1", x"0a53", x"08bb", x"0482", 
            x"feb6", x"fa08", x"f8c7", x"fa8d", 
            x"fcb3", x"fd37", x"fca0", x"fc56", 
            x"fcd5", x"fd52", x"fcfc", x"fc1d", 
            x"fb03", x"f9bd", x"f8df", x"f920", 
            x"fab2", x"fd2d", x"ff8a", x"00c1", 
            x"00b2", x"0029", x"000e", x"0001", 
            x"ff24", x"fdcd", x"fd19", x"fd95", 
            x"feca", x"001d", x"01ad", x"0368", 
            x"04b2", x"0503", x"0478", x"0352", 
            x"0140", x"fdd6", x"f9bd", x"f6b7", 
            x"f5ab", x"f56e", x"f473", x"f2e1", 
            x"f1b8", x"f0b6", x"eee3", x"ec40", 
            x"e99c", x"e7ad", x"e705", x"e859", 
            x"eb9d", x"ef90", x"f294", x"f450", 
            x"f5c5", x"f7a7", x"f974", x"fa57", 
            x"fa2a", x"f963", x"f8bf", x"f8b8", 
            x"f8f0", x"f8f8", x"f93b", x"fa37", 
            x"fba1", x"fcd2", x"fd4d", x"fd35", 
            x"fd53", x"fe8e", x"0142", x"0432", 
            x"0570", x"04bc", x"03ab", x"0364", 
            x"032e", x"01aa", x"fefd", x"fcd7", 
            x"fc48", x"fcba", x"fd33", x"fdf2", 
            x"ffbe", x"0241", x"0439", x"0528", 
            x"058f", x"05cf", x"058a", x"0425", 
            x"01d2", x"ff5e", x"fd80", x"fcb8", 
            x"fced", x"fd30", x"fcf9", x"fcd3", 
            x"fdae", x"ff62", x"0094", x"0047", 
            x"fef9", x"fd82", x"fc57", x"fbd5", 
            x"fc99", x"feeb", x"01de", x"03a6", 
            x"03a2", x"0363", x"03fd", x"04a8", 
            x"049d", x"049a", x"05a0", x"076f", 
            x"08c5", x"0902", x"08a9", x"0848", 
            x"07bb", x"06e6", x"0614", x"0524", 
            x"0386", x"013a", x"ff0c", x"fd70", 
            x"fc2a", x"fae5", x"f9b6", x"f919", 
            x"f955", x"fa00", x"fa6a", x"fa30", 
            x"f990", x"f938", x"f99d", x"fa37", 
            x"fa23", x"f945", x"f89c", x"f8eb", 
            x"fa24", x"fc24", x"ff38", x"0367", 
            x"0755", x"0911", x"07ea", x"0525", 
            x"02bf", x"01e2", x"028a", x"03b9", 
            x"03f2", x"0292", x"0074", x"ff20", 
            x"ffa6", x"01f0", x"04ce", x"06de", 
            x"075c", x"06b0", x"05ef", x"0581", 
            x"0572", x"0620", x"07af", x"08d4", 
            x"075c", x"0309", x"fe71", x"fc4f", 
            x"fd57", x"0065", x"032d", x"03e8", 
            x"02c6", x"0122", x"ffe7", x"ff15", 
            x"fe7d", x"fe0a", x"fd8e", x"fccd", 
            x"fbe1", x"fb57", x"fbd1", x"fd62", 
            x"ff52", x"00ed", x"023d", x"03ac", 
            x"056b", x"0761", x"0940", x"0aac"
        ),
        -- Block 24
        (
            x"0b40", x"0acc", x"0a11", x"0a69", 
            x"0bdc", x"0cad", x"0b50", x"0835", 
            x"0544", x"03ab", x"02b6", x"013c", 
            x"ff7e", x"fef1", x"ffe7", x"00a8", 
            x"ff59", x"fc3a", x"f994", x"f8eb", 
            x"f958", x"f8fe", x"f77b", x"f600", 
            x"f59f", x"f698", x"f8b8", x"fbc6", 
            x"ff48", x"0274", x"048d", x"0592", 
            x"069f", x"0898", x"0aff", x"0cf0", 
            x"0e4e", x"0f2a", x"0f71", x"0f13", 
            x"0e40", x"0d94", x"0d7d", x"0d6a", 
            x"0c64", x"0a37", x"0778", x"04dc", 
            x"029e", x"0097", x"feaa", x"fce1", 
            x"fb00", x"f86b", x"f4e9", x"f15a", 
            x"eefd", x"ede2", x"ecdb", x"eb63", 
            x"ea71", x"eba5", x"ef88", x"f4ad", 
            x"f8df", x"fab0", x"fa88", x"fa17", 
            x"fa8e", x"fb68", x"fb20", x"f97e", 
            x"f808", x"f845", x"fa0e", x"fbf2", 
            x"fd39", x"fead", x"00ca", x"026a", 
            x"01fe", x"ffad", x"fd6a", x"fcdd", 
            x"fdcb", x"fee5", x"ff7f", x"ff9f", 
            x"ff16", x"fd95", x"fb7a", x"f967", 
            x"f78a", x"f604", x"f533", x"f50b", 
            x"f4f3", x"f48d", x"f45a", x"f51c", 
            x"f712", x"f9b2", x"fc1a", x"fe40", 
            x"0109", x"04d8", x"08c8", x"0b74", 
            x"0c7b", x"0cfd", x"0df4", x"0f03", 
            x"0f2e", x"0e40", x"0d19", x"0cc6", 
            x"0d1e", x"0cb3", x"0a82", x"0737", 
            x"04dd", x"0477", x"04b4", x"03a9", 
            x"0126", x"fee6", x"fe35", x"fe5f", 
            x"fdb3", x"fbac", x"f972", x"f891", 
            x"f9c1", x"fc6d", x"fefd", x"0026", 
            x"0008", x"ff81", x"feed", x"fe18", 
            x"fd49", x"fd51", x"fe44", x"ff5e", 
            x"002a", x"00d2", x"00f8", x"0038", 
            x"ff40", x"ff3b", x"0039", x"0186", 
            x"034f", x"0631", x"0969", x"0b26", 
            x"0aa8", x"092a", x"0827", x"07a8", 
            x"06b2", x"0479", x"01bf", x"00ae", 
            x"021f", x"0422", x"0401", x"01aa", 
            x"ff8d", x"ff71", x"007a", x"006c", 
            x"fe9a", x"fcea", x"fd00", x"fddc", 
            x"fd7a", x"fb96", x"f9d7", x"f9b5", 
            x"fb31", x"fdb0", x"0057", x"01a1", 
            x"00a1", x"fe1a", x"fb87", x"f9df", 
            x"f939", x"f933", x"f96f", x"f9e9", 
            x"fb41", x"fe0d", x"0137", x"02a5", 
            x"01a7", x"ff78", x"fd49", x"fafd", 
            x"f86c", x"f61c", x"f4f1", x"f559", 
            x"f73e", x"f9f9", x"fc66", x"fdb4", 
            x"fe0b", x"fe01", x"fdd1", x"fd52", 
            x"fcaf", x"fc7b", x"fcc2", x"fd05", 
            x"fcde", x"fc2c", x"fb40", x"fa61", 
            x"f98e", x"f8d6", x"f84b", x"f7eb", 
            x"f843", x"fa09", x"fd23", x"0074", 
            x"02a4", x"0371", x"03c3", x"0438", 
            x"048e", x"04a4", x"051f", x"0656", 
            x"0764", x"073a", x"05ab", x"0349", 
            x"00c3", x"fe7c", x"fc9a", x"fb1b", 
            x"f9fc", x"f9a9", x"fac5", x"fd2e", 
            x"ffc8", x"0175", x"01ec", x"01cb", 
            x"0179", x"0100", x"00a8", x"00ed", 
            x"01d1", x"026a", x"0218", x"011c", 
            x"0000", x"ff40", x"ffb0", x"019f", 
            x"042a", x"0626", x"0779", x"08cd", 
            x"0a63", x"0ba8", x"0c24", x"0bd8", 
            x"0ab0", x"08a8", x"06b3", x"062b", 
            x"0754", x"0963", x"0bab", x"0e3d", 
            x"10b0", x"11af", x"105d", x"0d14", 
            x"08e1", x"04c3", x"0108", x"fd97", 
            x"fade", x"f9a0", x"fa38", x"fbee", 
            x"fd4f", x"fd97", x"fd66", x"fdee", 
            x"ffbd", x"0242", x"049f", x"0679", 
            x"0785", x"073e", x"0569", x"02e9", 
            x"016d", x"0221", x"0461", x"0612", 
            x"0584", x"0329", x"0161", x"01db", 
            x"0441", x"06f0", x"0899", x"08a8", 
            x"0724", x"04f8", x"03be", x"0442", 
            x"0589", x"0594", x"034c", x"ffcc", 
            x"fd9e", x"fe63", x"00f5", x"02c4", 
            x"0288", x"00fe", x"ff61", x"fe43", 
            x"fda2", x"fd90", x"fdba", x"fce9", 
            x"faa0", x"f83a", x"f7a1", x"f93a", 
            x"fc25", x"ff8e", x"02be", x"04cb", 
            x"05c8", x"0682", x"06cc", x"056f", 
            x"0222", x"fe66", x"fc0b", x"fb9c", 
            x"fc4a", x"fd11", x"fd64", x"fd34", 
            x"fcf4", x"fd1a", x"fd74", x"fda9", 
            x"fe1a", x"feec", x"ff51", x"fea3", 
            x"fd85", x"fce8", x"fc71", x"fb35", 
            x"f944", x"f747", x"f56d", x"f354", 
            x"f118", x"efb5", x"f005", x"f1c6", 
            x"f40e", x"f5e1", x"f723", x"f8ba", 
            x"fb41", x"fdf4", x"ff81", x"ff6c", 
            x"fe27", x"fc42", x"fa24", x"f8a5", 
            x"f853", x"f8e2", x"f9b3", x"fab6", 
            x"fc24", x"fdce", x"ff8b", x"0120", 
            x"01dd", x"015e", x"0015", x"febc", 
            x"fd69", x"fb89", x"f93e", x"f801", 
            x"f910", x"fbd1", x"fe59", x"ff84", 
            x"ffd6", x"fff5", x"ff93", x"fdfb", 
            x"fb5b", x"f8bd", x"f70b", x"f6c5", 
            x"f843", x"faf7", x"fd1a", x"fd99", 
            x"fd9a", x"feb2", x"00be", x"02a3", 
            x"0425", x"05ad", x"0705", x"07c8", 
            x"0833", x"092b", x"0aee", x"0ce0", 
            x"0e34", x"0e3d", x"0c9c", x"0a0b", 
            x"0827", x"07df", x"08b2", x"095a", 
            x"091e", x"0856", x"07ef", x"0876", 
            x"09b8", x"0afe", x"0b99", x"0b58", 
            x"0a24", x"0814", x"05b7", x"03db", 
            x"02ff", x"0334", x"03d1", x"0384", 
            x"01ab", x"ff57", x"fe20", x"fe13", 
            x"fd72", x"fb6c", x"f958", x"f8de", 
            x"fa4e", x"fcd8", x"ff63", x"0112", 
            x"01ca", x"0262", x"03a3", x"0570", 
            x"0727", x"080e", x"07f4", x"0741", 
            x"065d", x"053a", x"0391", x"013b", 
            x"fe59", x"fbcc", x"faac", x"fb5d", 
            x"fcea", x"fdae", x"fcf3", x"fb23", 
            x"f88f", x"f52f", x"f154", x"ee3e", 
            x"ecee", x"ecb8", x"ec16", x"ea83", 
            x"e94b", x"ea26", x"ed10", x"efef", 
            x"f0bf", x"ef8f", x"ee1a", x"edfe", 
            x"efb9", x"f2f3", x"f6af", x"f98c", 
            x"fb2d", x"fc72", x"fe07", x"ffc5", 
            x"01af", x"0431", x"06e5", x"0866", 
            x"07f6", x"067f", x"054a", x"0494", 
            x"035e", x"00b0", x"fd2a", x"fad5", 
            x"faeb", x"fd05", x"ffc6", x"0197", 
            x"0186", x"ffa8", x"fcf4", x"fa88", 
            x"f956", x"f9d8", x"fb82", x"fd19", 
            x"fdef", x"fe36", x"fe9b", x"ff70", 
            x"0000", x"ffa4", x"ff16", x"0013", 
            x"0353", x"0731", x"0908", x"07eb", 
            x"051c", x"020d", x"ff17", x"fc6a", 
            x"fabf", x"fa66", x"fa85", x"fa5c", 
            x"faa9", x"fc2c", x"fe71", x"0087", 
            x"0211", x"02b4", x"021c", x"0107", 
            x"00ca", x"0196", x"022b", x"0147", 
            x"ff27", x"fd5c", x"fd54", x"fef1", 
            x"00ca", x"0157", x"ffe1", x"fda3", 
            x"fcc1", x"fdfe", x"005f", x"0296", 
            x"046d", x"0669", x"0857", x"0922", 
            x"0801", x"0571", x"035c", x"03bd", 
            x"05e2", x"06c3", x"049a", x"016a", 
            x"00b0", x"0307", x"05c6", x"0677", 
            x"0592", x"04e8", x"04cb", x"0412", 
            x"02fe", x"0350", x"0559", x"0712", 
            x"0688", x"0422", x"01f9", x"0168", 
            x"022e", x"03df", x"0656", x"0966", 
            x"0c91", x"0f1a", x"1021", x"0eaf", 
            x"0a8f", x"04d5", x"ff31", x"fb0f", 
            x"f8e8", x"f82e", x"f83b", x"f949", 
            x"fbf2", x"ff2b", x"00db", x"009d", 
            x"ffc6", x"ff2d", x"fe5c", x"fd37", 
            x"fcf2", x"fed0", x"0250", x"0581", 
            x"071a", x"07bc", x"08c7", x"0aa6", 
            x"0c3d", x"0c44", x"0a90", x"086e", 
            x"074b", x"0731", x"0727", x"0639", 
            x"0454", x"029e", x"021a", x"022b", 
            x"01a0", x"0060", x"ffa6", x"006c", 
            x"020b", x"0335", x"0386", x"039f", 
            x"03dc", x"03aa", x"027e", x"00b8", 
            x"ff67", x"feec", x"fe8f", x"fdfb", 
            x"fe55", x"00c0", x"04e2", x"08de", 
            x"0a84", x"0927", x"0680", x"052a", 
            x"05d4", x"06bb", x"062b", x"046d", 
            x"0290", x"00e1", x"ff6a", x"fec4", 
            x"ff20", x"ff35", x"fddd", x"fbc4", 
            x"fa76", x"faae", x"fbd3", x"fcdd", 
            x"fd2b", x"fcb0", x"fbff", x"fb59", 
            x"fa71", x"f8d1", x"f6bd", x"f55d", 
            x"f5b1", x"f77b", x"f9b6", x"fbc5", 
            x"fd99", x"ff76", x"0148", x"02ab", 
            x"03ec", x"0627", x"08de", x"0a0b", 
            x"092c", x"085d", x"097f", x"0b34", 
            x"0aa4", x"0771", x"03c0", x"0164", 
            x"008c", x"0040", x"0018", x"010d", 
            x"0377", x"05f5", x"0704", x"0688", 
            x"05a7", x"04c8", x"02b3", x"ff7a", 
            x"fdb3", x"ff9d", x"03a7", x"057f", 
            x"032f", x"ff80", x"fe89", x"00eb", 
            x"037d", x"03b3", x"029f", x"0270", 
            x"034b", x"03f8", x"0403", x"03b9", 
            x"02de", x"0130", x"ff63", x"fe3a", 
            x"fdbb", x"fd9c", x"fe6e", x"0131", 
            x"0504", x"06e8", x"04d7", x"0023", 
            x"fc39", x"fad3", x"fa47", x"f892", 
            x"f63c", x"f51f", x"f5a7", x"f696", 
            x"f732", x"f7da", x"f8aa", x"f937", 
            x"f980", x"f98a", x"f8cc", x"f6f4", 
            x"f496", x"f2c1", x"f1e5", x"f1aa", 
            x"f1f4", x"f303", x"f48b", x"f5c6", 
            x"f692", x"f7a2", x"f919", x"fa10", 
            x"f9d6", x"f947", x"f9bf", x"fb5c", 
            x"fce1", x"fcea", x"fb9d", x"fac6", 
            x"fb9d", x"fd56", x"fe82", x"ff0c", 
            x"004e", x"02f4", x"05ac", x"06a0", 
            x"055f", x"0343", x"01fb", x"01c1", 
            x"01c9", x"01b8", x"01dc", x"0274", 
            x"02c0", x"01b5", x"ff6d", x"fcc2", 
            x"fa4b", x"f827", x"f637", x"f4d6", 
            x"f4c3", x"f60d", x"f7bc", x"f8d6", 
            x"f91a", x"f8b5", x"f7df", x"f725", 
            x"f719", x"f7ad", x"f85e", x"f8fe", 
            x"f9b1", x"fa38", x"f9e6", x"f8d4", 
            x"f81b", x"f868", x"f965", x"faa0", 
            x"fc3d", x"fe1c", x"ff6c", x"ff7f", 
            x"febc", x"fdff", x"fdb4", x"fd8c", 
            x"fd12", x"fc40", x"fba9", x"fbe1", 
            x"fd46", x"0006", x"03b6", x"06d5", 
            x"07c3", x"0677", x"04c9", x"0489", 
            x"058b", x"060c", x"04ee", x"0250", 
            x"ff38", x"fd17", x"fc91", x"fd09", 
            x"fd6d", x"fd78", x"fda6", x"fe0a", 
            x"fe03", x"fd59", x"fd14", x"fe34", 
            x"fff6", x"0019", x"fdfe", x"fc46", 
            x"fdd4", x"0226", x"05df", x"067f", 
            x"0431", x"0115", x"ffbc", x"0114", 
            x"036e", x"0408", x"028a", x"01e8", 
            x"0465", x"0868", x"0aa7", x"09bf", 
            x"06d7", x"03a0", x"0110", x"ff52", 
            x"fe51", x"fe30", x"fed8", x"ff55", 
            x"fe95", x"fd1c", x"fca0", x"fd91", 
            x"fed6", x"0010", x"025e", x"061f", 
            x"09ac", x"0b4a", x"0b2d", x"0b25", 
            x"0c4f", x"0df0", x"0ecb", x"0e78", 
            x"0da2", x"0cf7", x"0c25", x"0ae6", 
            x"09e7", x"0a18", x"0b84", x"0ce6", 
            x"0d1c", x"0bf3", x"0a2b", x"08dc", 
            x"08c3", x"09dd", x"0af5", x"0aab", 
            x"08fb", x"0725", x"0657", x"06ae", 
            x"07a4", x"0893", x"0890", x"0718", 
            x"04d7", x"02a7", x"008a", x"fe2d", 
            x"fc3a", x"fbed", x"fd7f", x"ffff", 
            x"0228", x"034b", x"03ab", x"0427", 
            x"0515", x"05ed", x"05ba", x"03c2", 
            x"0071", x"fd56", x"fbb8", x"fb9f", 
            x"fbe9", x"fb4b", x"f9e3", x"f928", 
            x"fa1f", x"fc15", x"fd64", x"fd2b", 
            x"fbf6", x"fae1", x"fa8d", x"fabb", 
            x"fadc", x"fb18", x"fbe2", x"fd35", 
            x"fe79", x"ff4e", x"0018", x"0186", 
            x"03df", x"0688", x"080c", x"0724", 
            x"0473", x"0241", x"0243", x"040c", 
            x"05a2", x"0535", x"02e6", x"00a3", 
            x"0046", x"0229", x"0500", x"06b4", 
            x"0594", x"022f", x"ff05", x"fde5", 
            x"fde2", x"fc94", x"f956", x"f5ef", 
            x"f42c", x"f41f", x"f506", x"f6a3", 
            x"f895", x"f98d", x"f85a", x"f525", 
            x"f170", x"eee8", x"ee79", x"f000", 
            x"f2b0", x"f637", x"faa9", x"ff77"
        ),
        -- Block 23
        (
            x"02f6", x"03b9", x"01db", x"fec3", 
            x"fc18", x"fa9c", x"fa24", x"fa27", 
            x"fa10", x"f97b", x"f881", x"f7a4", 
            x"f708", x"f602", x"f421", x"f1d8", 
            x"f075", x"f114", x"f3d8", x"f795", 
            x"fa7d", x"fb63", x"fa4f", x"f7e8", 
            x"f4d5", x"f1e2", x"f027", x"f072", 
            x"f261", x"f4dc", x"f763", x"fa52", 
            x"fe32", x"02e4", x"0769", x"0a63", 
            x"0b03", x"098f", x"070a", x"0449", 
            x"01a2", x"ff8f", x"ff1a", x"00aa", 
            x"02fa", x"0466", x"0498", x"044b", 
            x"03f1", x"0326", x"0186", x"ffaa", 
            x"fea1", x"febe", x"ff3e", x"ff54", 
            x"ff07", x"fefd", x"ff55", x"ff5f", 
            x"fed0", x"fe5b", x"fecc", x"002c", 
            x"01ed", x"0344", x"03ce", x"0389", 
            x"029d", x"0127", x"ff2c", x"fcf1", 
            x"fb4f", x"fb0c", x"fc0a", x"fdd7", 
            x"004d", x"0331", x"0531", x"047c", 
            x"011b", x"fd16", x"fa3c", x"f913", 
            x"f9a8", x"fba7", x"fe35", x"0080", 
            x"024e", x"045a", x"070b", x"0991", 
            x"0acc", x"0a79", x"0946", x"07c7", 
            x"0660", x"05fc", x"075f", x"09de", 
            x"0bb4", x"0bbe", x"0ab5", x"098e", 
            x"07f9", x"0548", x"01bc", x"fe74", 
            x"fc9d", x"fc96", x"fdba", x"fe79", 
            x"fd79", x"fbb3", x"fb54", x"fc37", 
            x"fbe4", x"f93c", x"f5d5", x"f3af", 
            x"f370", x"f4f0", x"f7e7", x"fb7f", 
            x"fea1", x"00fb", x"0298", x"03a7", 
            x"048a", x"057e", x"0649", x"06b7", 
            x"0700", x"0778", x"07df", x"0772", 
            x"0666", x"05cf", x"05fc", x"05c5", 
            x"0416", x"0132", x"fe57", x"fc62", 
            x"fb65", x"fb3e", x"fbce", x"fcac", 
            x"fcf0", x"fbb8", x"f9b5", x"f8a3", 
            x"f8f1", x"f927", x"f848", x"f771", 
            x"f82a", x"f9f4", x"fae6", x"fa76", 
            x"fa84", x"fd02", x"0130", x"0443", 
            x"0469", x"026b", x"0091", x"0066", 
            x"013f", x"014c", x"ff9c", x"fd0a", 
            x"fb1d", x"fa97", x"fb7c", x"fd9e", 
            x"0054", x"025e", x"02f6", x"0284", 
            x"01b9", x"005d", x"fe1e", x"fbcf", 
            x"fac0", x"fb10", x"fbe1", x"fd13", 
            x"ff78", x"038b", x"07ee", x"0a35", 
            x"09b6", x"0812", x"06dd", x"0655", 
            x"05f8", x"0598", x"0542", x"04da", 
            x"0432", x"031a", x"0161", x"ff79", 
            x"feb1", x"ffb9", x"0141", x"017c", 
            x"004c", x"ff55", x"0029", x"0288", 
            x"04bc", x"0547", x"046d", x"03e8", 
            x"04f4", x"06fa", x"0908", x"0b09", 
            x"0cad", x"0d7c", x"0dfc", x"0f5d", 
            x"119f", x"137e", x"1463", x"14e0", 
            x"1522", x"1494", x"12d3", x"0ffd", 
            x"0cc3", x"0a18", x"0891", x"076f", 
            x"04ad", x"ffa4", x"faa3", x"f829", 
            x"f7ba", x"f6d8", x"f457", x"f1da", 
            x"f1e1", x"f4f1", x"f964", x"fd73", 
            x"0095", x"0310", x"050f", x"0679", 
            x"072a", x"079c", x"08a5", x"0ad7", 
            x"0dbe", x"1047", x"11ef", x"133f", 
            x"146f", x"1450", x"1230", x"0f4c", 
            x"0d10", x"0bac", x"0a9f", x"0a19", 
            x"0a9b", x"0b53", x"0a37", x"05b0", 
            x"fe9b", x"f7d3", x"f3de", x"f2cc", 
            x"f2a7", x"f236", x"f276", x"f491", 
            x"f7fd", x"fb7b", x"fe58", x"ffe4", 
            x"fedf", x"fb56", x"f7c0", x"f6f2", 
            x"f968", x"fcf7", x"ff7f", x"00cd", 
            x"0197", x"0230", x"02a7", x"0380", 
            x"0569", x"0805", x"095d", x"086a", 
            x"0694", x"0591", x"0506", x"0395", 
            x"012c", x"fe60", x"fb21", x"f7ce", 
            x"f5ab", x"f58d", x"f6fe", x"f8a9", 
            x"f9a6", x"fa15", x"fa64", x"fa99", 
            x"fa62", x"fa0a", x"fa7a", x"fbb5", 
            x"fca7", x"fcc4", x"fd07", x"fe33", 
            x"ff4f", x"ff11", x"fdfe", x"fdbd", 
            x"fed3", x"0021", x"009b", x"0047", 
            x"ffa6", x"ff0e", x"fe73", x"fde1", 
            x"fdd1", x"fe87", x"ff8f", x"0007", 
            x"ff60", x"fdc8", x"fbd4", x"fa30", 
            x"f9eb", x"fb12", x"fbd9", x"fa5d", 
            x"f721", x"f4ee", x"f5bf", x"f824", 
            x"f8ff", x"f722", x"f49f", x"f467", 
            x"f6e5", x"f9a0", x"fa3d", x"f888", 
            x"f633", x"f51c", x"f5b9", x"f742", 
            x"f8dc", x"fa48", x"fb98", x"fcf8", 
            x"fe6f", x"ffd9", x"00fb", x"015d", 
            x"00cb", x"0011", x"007e", x"0217", 
            x"033f", x"0256", x"ff7d", x"fcdf", 
            x"fc89", x"fdf2", x"fe93", x"fd27", 
            x"fad4", x"f9bc", x"fabf", x"fca4", 
            x"fd8b", x"fcb2", x"fabe", x"f924", 
            x"f90a", x"fa07", x"fa12", x"f80e", 
            x"f57b", x"f4bb", x"f698", x"f9ac", 
            x"fc33", x"fe32", x"0098", x"031b", 
            x"043a", x"0389", x"022e", x"0170", 
            x"0181", x"01aa", x"0112", x"ffa4", 
            x"fe29", x"fd53", x"fd2b", x"fd15", 
            x"fc75", x"fae3", x"f888", x"f66e", 
            x"f5d4", x"f69c", x"f773", x"f775", 
            x"f707", x"f6f0", x"f744", x"f7d6", 
            x"f890", x"f8b0", x"f713", x"f406", 
            x"f1c7", x"f23a", x"f4f4", x"f833", 
            x"fb14", x"fdb9", x"0076", x"0392", 
            x"06fe", x"09d7", x"0aef", x"0a49", 
            x"091d", x"0833", x"0720", x"0574", 
            x"03a3", x"025b", x"01c6", x"020a", 
            x"02ed", x"038e", x"031c", x"01b7", 
            x"001a", x"fef2", x"feab", x"ff3c", 
            x"ff76", x"fe22", x"fbda", x"fa7b", 
            x"faf7", x"fc88", x"fe04", x"feb0", 
            x"feb0", x"feb4", x"ff39", x"0065", 
            x"026a", x"04ef", x"06b7", x"0669", 
            x"03cf", x"0063", x"fdfd", x"fd4e", 
            x"fe2c", x"0000", x"0198", x"01f8", 
            x"015c", x"00e3", x"013c", x"0201", 
            x"0243", x"0182", x"0001", x"fe95", 
            x"fded", x"fde8", x"fe1c", x"fe88", 
            x"ff5a", x"0026", x"0018", x"fed3", 
            x"fcf4", x"fbc6", x"fc5b", x"fe7c", 
            x"0091", x"0127", x"00a3", x"00b4", 
            x"01c1", x"02e2", x"0362", x"02d3", 
            x"0124", x"ff7f", x"ff6c", x"014d", 
            x"03b9", x"04bc", x"035b", x"0018", 
            x"fca0", x"faa2", x"fa78", x"fb10", 
            x"fafc", x"f9c4", x"f8bb", x"f965", 
            x"fbb2", x"fe6e", x"0082", x"019e", 
            x"01db", x"01b7", x"01ec", x"02c1", 
            x"03cc", x"046e", x"04d5", x"05cc", 
            x"077c", x"090f", x"09a5", x"0960", 
            x"0901", x"08bd", x"07ba", x"04ca", 
            x"003a", x"fcc8", x"fd32", x"009a", 
            x"0350", x"033d", x"0191", x"fffb", 
            x"fe61", x"fc34", x"fa6b", x"fa6f", 
            x"fc3d", x"fe72", x"ff92", x"ff80", 
            x"ff6e", x"0071", x"0292", x"04a5", 
            x"057b", x"0547", x"04d2", x"0413", 
            x"02cf", x"01e3", x"02c7", x"05ac", 
            x"08b2", x"09b9", x"08e9", x"0885", 
            x"0a29", x"0cc8", x"0e0f", x"0cdb", 
            x"097d", x"04c9", x"ffc2", x"fbc5", 
            x"fa0c", x"fad9", x"fd56", x"000f", 
            x"01c9", x"0246", x"027c", x"0372", 
            x"0478", x"03c2", x"0104", x"fdef", 
            x"fc38", x"fb8c", x"fa2c", x"f7c1", 
            x"f64f", x"f7c7", x"fb7a", x"fe89", 
            x"ff36", x"fe6b", x"fe57", x"0018", 
            x"02d3", x"04f2", x"0551", x"03be", 
            x"00e9", x"fe83", x"fe5d", x"00d1", 
            x"040d", x"0588", x"04ae", x"0374", 
            x"03fa", x"05f2", x"0769", x"0727", 
            x"0612", x"0592", x"059e", x"059e", 
            x"05b9", x"0651", x"0714", x"0726", 
            x"05ce", x"037c", x"01cb", x"019a", 
            x"01d5", x"00be", x"fdea", x"fae3", 
            x"f962", x"f96e", x"f9b3", x"f9a2", 
            x"f9fa", x"fb63", x"fd51", x"feaa", 
            x"fee0", x"fe8f", x"fed0", x"ffe9", 
            x"00ec", x"00bf", x"ff38", x"fdc7", 
            x"fe57", x"00f5", x"03b5", x"0525", 
            x"05a5", x"0630", x"0714", x"07dd", 
            x"0802", x"07b0", x"0771", x"0754", 
            x"0705", x"05b7", x"0352", x"017d", 
            x"01f0", x"043e", x"0626", x"05cf", 
            x"03eb", x"02f5", x"03ba", x"04c1", 
            x"047f", x"02f3", x"016b", x"014e", 
            x"0316", x"05c4", x"07ac", x"0845", 
            x"0870", x"0892", x"0850", x"0757", 
            x"0588", x"0270", x"fdd8", x"f92a", 
            x"f6c4", x"f753", x"f9b4", x"fd20", 
            x"0142", x"0501", x"06a7", x"05a9", 
            x"031f", x"006f", x"fe20", x"fc4c", 
            x"faec", x"f9b4", x"f8b5", x"f89e", 
            x"f978", x"fa24", x"fa09", x"fa2e", 
            x"fb86", x"fd61", x"fe6a", x"fe76", 
            x"fe02", x"fce6", x"fb0d", x"f95c", 
            x"f96e", x"fb8a", x"fdb2", x"fde0", 
            x"fc78", x"fba1", x"fc86", x"fe5b", 
            x"ffd3", x"0064", x"0091", x"0131", 
            x"02cc", x"0524", x"0750", x"0815", 
            x"06ea", x"049e", x"025b", x"00da", 
            x"008b", x"0101", x"00e7", x"ffa9", 
            x"fe74", x"fef2", x"00a9", x"0188", 
            x"00fe", x"00b0", x"018b", x"01fe", 
            x"00e4", x"ff5f", x"feea", x"ff2a", 
            x"ff15", x"ff29", x"006d", x"0241", 
            x"031d", x"029d", x"0192", x"00a0", 
            x"ffde", x"ff57", x"ff38", x"ff4f", 
            x"fefd", x"fd7a", x"faf8", x"f8fe", 
            x"f90f", x"fae3", x"fc37", x"fb6e", 
            x"f977", x"f832", x"f816", x"f833", 
            x"f80f", x"f865", x"f9ae", x"fb31", 
            x"fbde", x"fbad", x"fbc4", x"fd6d", 
            x"00dc", x"04e1", x"07f9", x"0986", 
            x"09ed", x"09e6", x"09ee", x"0a16", 
            x"0a02", x"091f", x"0772", x"055c", 
            x"02e9", x"0037", x"fe01", x"fd84", 
            x"fefb", x"009a", x"0034", x"fd82", 
            x"fa76", x"f8e0", x"f893", x"f83d", 
            x"f705", x"f4f9", x"f2c4", x"f0f9", 
            x"ef52", x"ed41", x"eb5c", x"eb54", 
            x"ed9a", x"f033", x"f115", x"f0c9", 
            x"f142", x"f31c", x"f564", x"f777", 
            x"f931", x"fa08", x"f9c4", x"f9e5", 
            x"fc8a", x"0161", x"062f", x"0985", 
            x"0b9c", x"0cbf", x"0ca5", x"0b3f", 
            x"0944", x"07b9", x"0709", x"0647", 
            x"043a", x"0181", x"003b", x"0161", 
            x"03a1", x"0531", x"0586", x"0528", 
            x"0488", x"03c6", x"031b", x"0271", 
            x"0184", x"00ab", x"0031", x"ffa1", 
            x"fe8a", x"fde0", x"fec5", x"00dd", 
            x"02e0", x"0430", x"04ec", x"050f", 
            x"048b", x"0396", x"026b", x"00b9", 
            x"fe35", x"fb77", x"f9e7", x"fa9a", 
            x"fd02", x"ffa6", x"0139", x"0130", 
            x"ffd8", x"fe33", x"fd56", x"fdd2", 
            x"ff11", x"ff7f", x"fe5d", x"fd28", 
            x"fdce", x"ffbc", x"0073", x"fe7f", 
            x"faf6", x"f856", x"f827", x"f9ef", 
            x"fc5d", x"ff23", x"02aa", x"061a", 
            x"06e4", x"03c2", x"ff13", x"fc2f", 
            x"fc23", x"fd4a", x"fdd3", x"fdda", 
            x"fee0", x"01b5", x"05a0", x"0912", 
            x"0ab0", x"0a50", x"08df", x"0747", 
            x"05bc", x"0441", x"030f", x"0243", 
            x"01be", x"0194", x"020b", x"0318", 
            x"0420", x"03c8", x"00f1", x"fc6d", 
            x"f91a", x"f8df", x"fa52", x"fac8", 
            x"fa51", x"fb54", x"fe25", x"0038", 
            x"ffe2", x"feb8", x"ff0e", x"0089", 
            x"00ae", x"fe9d", x"fc06", x"fb4c", 
            x"fd58", x"0072", x"01c1", x"0024", 
            x"fd4c", x"fbe9", x"fcf2", x"ff11", 
            x"00e1", x"0224", x"02cb", x"0241", 
            x"001e", x"fd0f", x"fa98", x"f981", 
            x"f95a", x"f9f5", x"fc43", x"010d", 
            x"06b3", x"09ed", x"0983", x"079c", 
            x"06c3", x"0742", x"07e3", x"07ad", 
            x"068f", x"052c", x"0446", x"048f", 
            x"0648", x"08b7", x"0a44", x"09ae", 
            x"0776", x"055b", x"0466", x"039a", 
            x"0184", x"fe2a", x"fb29", x"fa03", 
            x"fa46", x"fa54", x"f9aa", x"f961", 
            x"fac7", x"fd74", x"ff4b", x"feec", 
            x"fd16", x"fb58", x"fa79", x"fa9f", 
            x"fbc4", x"fda1", x"ff61", x"003c", 
            x"008b", x"01c2", x"04a2", x"0846", 
            x"0aec", x"0b3f", x"097c", x"0736", 
            x"0581", x"03e0", x"0229", x"01fd"
        ),
        -- Block 22
        (
            x"049b", x"083b", x"09ea", x"0982", 
            x"095c", x"0a77", x"0b32", x"09f9", 
            x"0787", x"057b", x"0405", x"01ff", 
            x"ff28", x"fd8a", x"ff59", x"039f", 
            x"0665", x"0524", x"01cb", x"fff7", 
            x"0052", x"0086", x"ff15", x"fd27", 
            x"fcaa", x"fe38", x"00ef", x"034c", 
            x"03db", x"02be", x"01c6", x"0186", 
            x"000e", x"fba8", x"f5bd", x"f241", 
            x"f3d3", x"f83b", x"fa94", x"f8fa", 
            x"f616", x"f575", x"f756", x"f94f", 
            x"f9e6", x"fa24", x"fba2", x"fea8", 
            x"0216", x"040d", x"0345", x"0081", 
            x"fd9a", x"fb8b", x"fa5f", x"fa4d", 
            x"fbd3", x"fe66", x"00c2", x"0241", 
            x"02d4", x"0259", x"0089", x"fdda", 
            x"fbc3", x"fb78", x"fcab", x"fdd4", 
            x"fdc9", x"fcc3", x"fba8", x"fab1", 
            x"f9b2", x"f89f", x"f746", x"f575", 
            x"f3a8", x"f2aa", x"f324", x"f51e", 
            x"f77b", x"f8a2", x"f7b2", x"f4f0", 
            x"f158", x"ee75", x"ed9b", x"eeff", 
            x"f18c", x"f334", x"f30d", x"f2c9", 
            x"f49c", x"f812", x"fa7e", x"fa20", 
            x"f7bf", x"f4ef", x"f2a5", x"f18e", 
            x"f1b9", x"f2ad", x"f3f9", x"f571", 
            x"f719", x"f8cd", x"fa52", x"fbb4", 
            x"fd28", x"ff1a", x"01d5", x"048f", 
            x"0565", x"03d2", x"0225", x"02c9", 
            x"04f5", x"05cf", x"0427", x"0148", 
            x"ff8c", x"0076", x"0344", x"0579", 
            x"0585", x"0404", x"026b", x"00f2", 
            x"ff41", x"fe14", x"fe4e", x"ff4d", 
            x"ffa5", x"ff06", x"fe1c", x"fd53", 
            x"fc98", x"fbc4", x"facc", x"fa72", 
            x"fc07", x"ff8a", x"02a6", x"0381", 
            x"038a", x"0573", x"0929", x"0be1", 
            x"0bee", x"0ac3", x"0a65", x"0a4b", 
            x"08fb", x"0660", x"03e8", x"0352", 
            x"052c", x"07c1", x"08ce", x"0847", 
            x"0846", x"09fe", x"0c21", x"0d17", 
            x"0cdf", x"0d06", x"0e7c", x"0fe5", 
            x"0f90", x"0e1e", x"0d90", x"0ebf", 
            x"10cf", x"121e", x"1197", x"0f75", 
            x"0cee", x"0b17", x"09fd", x"087c", 
            x"05de", x"035f", x"02c5", x"03db", 
            x"047f", x"038a", x"01db", x"007d", 
            x"ff45", x"fd92", x"fb6b", x"f994", 
            x"f88a", x"f870", x"f99e", x"fc3b", 
            x"ff5d", x"016d", x"01cf", x"0146", 
            x"00d1", x"0062", x"0028", x"015e", 
            x"0495", x"083a", x"09c6", x"08a7", 
            x"06e1", x"06de", x"091c", x"0bbf", 
            x"0c39", x"0a03", x"0748", x"063e", 
            x"06b7", x"0665", x"03d4", x"002e", 
            x"fde3", x"fdd4", x"fe87", x"fe8a", 
            x"fe44", x"fe89", x"febe", x"fd8f", 
            x"fb22", x"f984", x"fa27", x"fbc7", 
            x"fc9e", x"fd07", x"fea1", x"0116", 
            x"0290", x"02c9", x"0355", x"0514", 
            x"06f7", x"07c6", x"079f", x"06f5", 
            x"05b5", x"0438", x"03bc", x"04bd", 
            x"05db", x"05e8", x"0550", x"04ad", 
            x"0351", x"00cc", x"fde4", x"fb61", 
            x"f980", x"f86b", x"f878", x"f9d9", 
            x"fcc5", x"0126", x"064c", x"09ed", 
            x"0927", x"0416", x"fe9a", x"fc9a", 
            x"fdd6", x"ff39", x"ffab", x"00ff", 
            x"0487", x"08be", x"0b02", x"0a66", 
            x"07e0", x"04df", x"01eb", x"febb", 
            x"faea", x"f73c", x"f628", x"f92d", 
            x"fe93", x"029a", x"0369", x"0267", 
            x"0106", x"fea4", x"faa9", x"f70f", 
            x"f60f", x"f6ef", x"f728", x"f5f1", 
            x"f4d5", x"f531", x"f6b9", x"f826", 
            x"f7fb", x"f551", x"f14a", x"eeb4", 
            x"ef90", x"f327", x"f6f5", x"f94c", 
            x"fa46", x"faef", x"fba9", x"fbd3", 
            x"facb", x"f95c", x"f936", x"fa99", 
            x"fbc2", x"fb48", x"fa0e", x"f9b2", 
            x"fa4b", x"fb23", x"fc50", x"fe45", 
            x"003d", x"00ac", x"fef5", x"fbbb", 
            x"f889", x"f707", x"f7d0", x"f9bd", 
            x"faa0", x"f96c", x"f7a9", x"f7b6", 
            x"fa29", x"fd33", x"fe4c", x"fcf1", 
            x"fb4b", x"fbe1", x"ff11", x"02e0", 
            x"0534", x"05b9", x"0539", x"04ba", 
            x"04dd", x"0590", x"066a", x"0786", 
            x"093b", x"0adb", x"0b0b", x"09b5", 
            x"085b", x"07d3", x"0752", x"0635", 
            x"04e7", x"0380", x"0150", x"fe51", 
            x"fb79", x"f9d1", x"f9b1", x"fab3", 
            x"fbd4", x"fbd3", x"fa52", x"f8a4", 
            x"f81e", x"f8ab", x"f929", x"f8b8", 
            x"f7f6", x"f8a8", x"fbf3", x"00bf", 
            x"0473", x"05fa", x"06a2", x"07db", 
            x"0911", x"08ee", x"07bd", x"06a0", 
            x"0628", x"06a1", x"081a", x"099f", 
            x"09e0", x"0909", x"087b", x"08d0", 
            x"08e9", x"078b", x"04ce", x"012b", 
            x"fccf", x"f90f", x"f875", x"fb37", 
            x"fde3", x"fdaf", x"fbdd", x"faf6", 
            x"fab1", x"f916", x"f66d", x"f536", 
            x"f6a2", x"f949", x"fb6d", x"fc87", 
            x"fc88", x"fb59", x"fa1b", x"fb2d", 
            x"ffbd", x"05a3", x"0928", x"099d", 
            x"0a78", x"0ef9", x"15d3", x"1a52", 
            x"19ac", x"156b", x"1086", x"0bf7", 
            x"0758", x"0311", x"00b9", x"00cd", 
            x"01b0", x"0253", x"03a5", x"0650", 
            x"0899", x"0782", x"027c", x"fc5f", 
            x"f831", x"f75d", x"f9d2", x"fe02", 
            x"01c3", x"043a", x"059f", x"05a4", 
            x"036b", x"ffbc", x"fd9a", x"fea5", 
            x"00fa", x"01d4", x"0131", x"0145", 
            x"0336", x"05da", x"07a3", x"088d", 
            x"0890", x"0693", x"0269", x"fe7f", 
            x"fd90", x"ff85", x"01fc", x"02ff", 
            x"0225", x"ffda", x"fd2c", x"fb56", 
            x"fad5", x"fabf", x"f9bc", x"f785", 
            x"f58d", x"f4ef", x"f549", x"f5da", 
            x"f620", x"f5d0", x"f50a", x"f433", 
            x"f3b2", x"f466", x"f73e", x"fb58", 
            x"fdcd", x"fc89", x"f92f", x"f72a", 
            x"f7c6", x"f97d", x"fa52", x"f9a5", 
            x"f845", x"f812", x"fa80", x"fe92", 
            x"0141", x"007d", x"fd90", x"fba8", 
            x"fcfe", x"011e", x"055f", x"074a", 
            x"0664", x"041b", x"01c4", x"ffec", 
            x"fef9", x"ff04", x"ff08", x"fdce", 
            x"fb92", x"fa07", x"fa17", x"fb0a", 
            x"fbd5", x"fc3f", x"fc47", x"fb42", 
            x"f8fd", x"f67c", x"f529", x"f56e", 
            x"f631", x"f5f2", x"f473", x"f2cf", 
            x"f254", x"f3a1", x"f665", x"f977", 
            x"fb80", x"fbbd", x"fac6", x"f9ff", 
            x"fa5b", x"fb7b", x"fc78", x"fcf6", 
            x"fd84", x"feb1", x"ffee", x"012e", 
            x"03ac", x"0791", x"0a3a", x"08b6", 
            x"03c7", x"ff58", x"fe01", x"fe94", 
            x"fe93", x"fd6f", x"fc8a", x"fcfa", 
            x"fe51", x"fefb", x"fd42", x"f8dd", 
            x"f383", x"ef4f", x"ed5d", x"eda6", 
            x"ef7f", x"f1f9", x"f402", x"f50a", 
            x"f561", x"f60d", x"f7c1", x"fa17", 
            x"fc16", x"fd56", x"fe1b", x"fee4", 
            x"0062", x"038e", x"0886", x"0dca", 
            x"11ad", x"1475", x"17b1", x"1b65", 
            x"1d2b", x"1b95", x"1877", x"15d5", 
            x"12c5", x"0e22", x"0a26", x"09db", 
            x"0c9c", x"0ec0", x"0df2", x"0b01", 
            x"0812", x"0668", x"05bf", x"04ae", 
            x"021c", x"fe40", x"fa82", x"f878", 
            x"f841", x"f89a", x"f8d5", x"f996", 
            x"fc04", x"0054", x"04ba", x"078e", 
            x"096a", x"0b5f", x"0d05", x"0d9e", 
            x"0de5", x"0f10", x"10fc", x"12c3", 
            x"13b7", x"136d", x"11fa", x"0ff7", 
            x"0dad", x"0b22", x"0919", x"084b", 
            x"0798", x"053f", x"01d1", x"004c", 
            x"0291", x"06bf", x"09b1", x"0a32", 
            x"08fc", x"071c", x"0565", x"0456", 
            x"0381", x"01cf", x"ff53", x"fd49", 
            x"fc25", x"fb3e", x"fa5d", x"fa76", 
            x"fc47", x"ff08", x"0100", x"013b", 
            x"000b", x"fee9", x"ffac", x"0311", 
            x"072d", x"0858", x"0527", x"0071", 
            x"fe51", x"ff48", x"ffde", x"fd71", 
            x"f9fc", x"f9d3", x"fdca", x"01f7", 
            x"0256", x"fe99", x"f9d2", x"f769", 
            x"f84d", x"fa85", x"fb44", x"f9b8", 
            x"f83a", x"f9b8", x"fdfb", x"01e5", 
            x"0326", x"0253", x"017e", x"0182", 
            x"016b", x"0039", x"feaa", x"fe79", 
            x"0013", x"01f9", x"02b4", x"02be", 
            x"0328", x"038b", x"0348", x"02f0", 
            x"02a8", x"017a", x"ff2f", x"fd58", 
            x"fcec", x"fca6", x"fb31", x"f95b", 
            x"f898", x"f8ba", x"f851", x"f64d", 
            x"f310", x"efd7", x"edf5", x"edf7", 
            x"ef4a", x"f0cc", x"f228", x"f3a4", 
            x"f4c1", x"f497", x"f2f9", x"f112", 
            x"f12f", x"f4ba", x"fa67", x"fe8c", 
            x"fe9b", x"fc61", x"fc0e", x"ff6c", 
            x"042d", x"06ed", x"069a", x"050b", 
            x"049f", x"05b8", x"072d", x"0830", 
            x"0889", x"07ab", x"058d", x"0363", 
            x"01b0", x"ff8e", x"fcba", x"fab9", 
            x"fa98", x"fb9b", x"fd3d", x"fff9", 
            x"0316", x"044e", x"02c3", x"0090", 
            x"0015", x"009e", x"ff7f", x"fc07", 
            x"f8bb", x"f83e", x"fa76", x"fcf9", 
            x"fe02", x"fdf3", x"fe19", x"fe99", 
            x"fec6", x"febd", x"ff27", x"0017", 
            x"01a0", x"0429", x"06d0", x"075a", 
            x"04e2", x"0134", x"fe49", x"fc5c", 
            x"fab3", x"f92f", x"f7e0", x"f64c", 
            x"f46f", x"f327", x"f32a", x"f46a", 
            x"f6a4", x"f92b", x"fac2", x"fa8f", 
            x"f906", x"f800", x"f943", x"fc22", 
            x"fdf7", x"fd5d", x"fbdc", x"fb98", 
            x"fc53", x"fc56", x"fbaa", x"fc69", 
            x"ffbc", x"03dd", x"0635", x"06b2", 
            x"076d", x"0973", x"0ae3", x"092f", 
            x"04bd", x"00a5", x"ff0f", x"ff82", 
            x"00a4", x"017e", x"0160", x"003c", 
            x"ff14", x"fede", x"ff7a", x"002a", 
            x"0073", x"0037", x"ff52", x"fe6a", 
            x"fefd", x"0104", x"0229", x"0100", 
            x"fe92", x"fc78", x"fb1e", x"fa72", 
            x"fb2d", x"fd8b", x"0021", x"0157", 
            x"0167", x"019b", x"0229", x"0282", 
            x"0326", x"04ff", x"0762", x"0888", 
            x"081e", x"0784", x"07b0", x"0842", 
            x"08d8", x"09af", x"0ab6", x"0afe", 
            x"0a33", x"097d", x"09d4", x"0a47", 
            x"097f", x"082f", x"07c0", x"082b", 
            x"087c", x"0823", x"0747", x"066b", 
            x"060e", x"06bc", x"0824", x"08d9", 
            x"0822", x"06b5", x"05a3", x"0553", 
            x"0532", x"0437", x"0201", x"ff4a", 
            x"fd0d", x"fc16", x"fcf5", x"ffc6", 
            x"03b7", x"06e6", x"076f", x"04d2", 
            x"0032", x"fbd7", x"f9cf", x"fa9b", 
            x"fceb", x"ff34", x"0086", x"0073", 
            x"ff87", x"ff50", x"007b", x"015a", 
            x"fff7", x"fce3", x"fa74", x"fa32", 
            x"fbae", x"fd92", x"fea2", x"febc", 
            x"fedd", x"ff77", x"ff92", x"fe8a", 
            x"fdf2", x"0029", x"04a2", x"0821", 
            x"0906", x"08fd", x"0a79", x"0d94", 
            x"0fdf", x"0f7d", x"0d54", x"0b83", 
            x"0ad3", x"09fa", x"073b", x"02c0", 
            x"fec1", x"fccd", x"fcb7", x"fce9", 
            x"fbd5", x"f960", x"f6eb", x"f608", 
            x"f748", x"fa26", x"fdb0", x"009d", 
            x"00fb", x"fe3f", x"fb24", x"fad7", 
            x"fc49", x"fb42", x"f673", x"f201", 
            x"f28c", x"f78f", x"fc89", x"fea6", 
            x"feec", x"fefd", x"feb0", x"fd78", 
            x"fbd2", x"fa27", x"f7d6", x"f528", 
            x"f4aa", x"f82f", x"fd3a", x"feec", 
            x"fbbf", x"f794", x"f6d0", x"f9d1", 
            x"fe0e", x"011a", x"0191", x"ff45", 
            x"fb77", x"f7db", x"f49f", x"f09c", 
            x"eb98", x"e77e", x"e6bb", x"e9f7", 
            x"ef63", x"f3fc", x"f64c", x"f76d", 
            x"f919", x"fb60", x"fd5c", x"ff12", 
            x"00ea", x"02bd", x"04ab", x"0754", 
            x"0a37", x"0b7b", x"0a4f", x"080b", 
            x"063d", x"04b7", x"0348", x"0310", 
            x"042e", x"04c4", x"038f", x"01d3", 
            x"009a", x"fdf7", x"f82b", x"f18f", 
            x"ee56", x"ef95", x"f225", x"f209", 
            x"ee9f", x"eaa4", x"e8f5", x"ea35", 
            x"eccc", x"eec4", x"efae", x"f0e6"
        ),
        -- Block 21
        (
            x"f3f7", x"f888", x"fc6a", x"fe03", 
            x"fdaa", x"fcb8", x"fc00", x"fb2d", 
            x"f9b7", x"f7f6", x"f781", x"fa38", 
            x"ffba", x"04cc", x"06f5", x"0779", 
            x"09ad", x"0f46", x"159b", x"1739", 
            x"1237", x"0b1d", x"07fa", x"09f3", 
            x"0d28", x"0da8", x"0b2f", x"0860", 
            x"076c", x"0818", x"0845", x"060a", 
            x"01ca", x"fde8", x"fc04", x"fb84", 
            x"faf8", x"fa15", x"f98e", x"f9ed", 
            x"fa89", x"f9f7", x"f7b6", x"f5a8", 
            x"f67e", x"fa1a", x"fd2b", x"fd81", 
            x"fc5e", x"fc39", x"fdb6", x"ffbd", 
            x"017c", x"0316", x"048d", x"04dd", 
            x"0365", x"01ec", x"02e3", x"060c", 
            x"08a4", x"08ce", x"07a1", x"069d", 
            x"0543", x"0340", x"0260", x"03c7", 
            x"05ea", x"06cf", x"064f", x"0534", 
            x"0406", x"03fa", x"0685", x"0a9b", 
            x"0d4d", x"0d5b", x"0bd9", x"09e3", 
            x"088a", x"0952", x"0c2d", x"0e19", 
            x"0cbf", x"09c5", x"0840", x"0895", 
            x"0946", x"0984", x"093e", x"08c0", 
            x"08e6", x"0a5b", x"0ba9", x"0a5d", 
            x"06ed", x"0456", x"03b5", x"02f7", 
            x"00a4", x"fe65", x"fe98", x"00be", 
            x"0216", x"014c", x"0011", x"0020", 
            x"0090", x"ff6e", x"fcf2", x"fb93", 
            x"fcee", x"ffbd", x"01ad", x"021f", 
            x"01cc", x"015f", x"0114", x"0122", 
            x"01b0", x"02ff", x"055f", x"0871", 
            x"0b06", x"0bcc", x"0a3a", x"06fb", 
            x"03e3", x"02ac", x"03a0", x"05ff", 
            x"08c3", x"0b68", x"0e43", x"11d8", 
            x"1501", x"15ab", x"12e5", x"0e18", 
            x"09b1", x"06cf", x"052a", x"0423", 
            x"034f", x"0260", x"014d", x"0035", 
            x"ff0b", x"fd56", x"fab2", x"f797", 
            x"f523", x"f369", x"f17e", x"ef2b", 
            x"ed2f", x"ec54", x"ed4c", x"f024", 
            x"f3dc", x"f720", x"f9ab", x"fc22", 
            x"fed5", x"019a", x"03ff", x"04ea", 
            x"03c7", x"0234", x"02bc", x"05ab", 
            x"077f", x"0501", x"0000", x"fd82", 
            x"ff91", x"032c", x"0415", x"01cf", 
            x"ffce", x"0046", x"0186", x"017d", 
            x"0156", x"036b", x"0710", x"087e", 
            x"0536", x"ff79", x"fbe8", x"fc77", 
            x"feb9", x"ff9a", x"ff05", x"fe9b", 
            x"fe98", x"fe02", x"fd91", x"ff74", 
            x"0414", x"089e", x"09d8", x"0713", 
            x"0267", x"ff4b", x"fffd", x"03be", 
            x"079f", x"094a", x"08c8", x"072f", 
            x"0531", x"03ec", x"048a", x"0652", 
            x"06b2", x"03f5", x"ff8b", x"fc5d", 
            x"fb9c", x"fbd7", x"faff", x"f8a3", 
            x"f604", x"f41e", x"f280", x"f066", 
            x"ee4e", x"edd3", x"efd6", x"f36a", 
            x"f6a9", x"f886", x"f94d", x"f986", 
            x"f971", x"f961", x"f985", x"f963", 
            x"f838", x"f647", x"f591", x"f833", 
            x"fdd2", x"0440", x"0976", x"0c0d", 
            x"0b6b", x"082f", x"040c", x"0072", 
            x"fdbe", x"fb97", x"f964", x"f6d0", 
            x"f4a7", x"f41c", x"f50c", x"f612", 
            x"f61f", x"f56a", x"f4e2", x"f434", 
            x"f20e", x"ee69", x"eb66", x"eb5e", 
            x"ee7e", x"f2be", x"f684", x"fa04", 
            x"fdc8", x"009f", x"00a7", x"fe35", 
            x"fbca", x"faf9", x"faef", x"faae", 
            x"fb11", x"fd3f", x"0048", x"0223", 
            x"024f", x"01d7", x"01b3", x"01c0", 
            x"0113", x"ff48", x"fd63", x"fc46", 
            x"fb4f", x"fa04", x"f9c8", x"fbf4", 
            x"fed4", x"ff4a", x"fd09", x"fb1d", 
            x"fb95", x"fd71", x"ffb4", x"0344", 
            x"081b", x"0b94", x"0bbf", x"09c8", 
            x"083c", x"083c", x"08b3", x"07e4", 
            x"05bf", x"0378", x"01cb", x"013b", 
            x"02bd", x"0661", x"0997", x"094b", 
            x"05c1", x"0256", x"0152", x"022b", 
            x"03b3", x"05bb", x"08a6", x"0c10", 
            x"0f1c", x"1114", x"11ab", x"10ed", 
            x"0f81", x"0e5a", x"0e2b", x"0ed3", 
            x"0ef3", x"0d29", x"09ad", x"0641", 
            x"041c", x"02c0", x"016b", x"0048", 
            x"fff3", x"001b", x"ffb6", x"fe46", 
            x"fc30", x"f9f1", x"f7e1", x"f65e", 
            x"f5c0", x"f648", x"f757", x"f76b", 
            x"f602", x"f4ca", x"f5f5", x"f9ed", 
            x"fe70", x"007f", x"ff30", x"fc4c", 
            x"fa77", x"fabd", x"fc47", x"fdf7", 
            x"ff2c", x"ff5a", x"fe91", x"fe85", 
            x"0131", x"0615", x"0a29", x"0aa8", 
            x"07c1", x"0468", x"0314", x"02ef", 
            x"0130", x"fd68", x"fa9f", x"fba9", 
            x"ff3e", x"015f", x"ffe5", x"fbfd", 
            x"f84a", x"f6a5", x"f705", x"f7db", 
            x"f7eb", x"f7a9", x"f7b8", x"f773", 
            x"f694", x"f639", x"f74b", x"f8f3", 
            x"fa1c", x"fb1e", x"fc82", x"fe15", 
            x"fff1", x"02cb", x"0601", x"077c", 
            x"065d", x"041a", x"0272", x"01e2", 
            x"0186", x"000b", x"fd26", x"fa2d", 
            x"f8ca", x"f87f", x"f782", x"f58e", 
            x"f416", x"f3c7", x"f30a", x"f026", 
            x"ec59", x"ea73", x"eb89", x"ee58", 
            x"f101", x"f2cd", x"f4cc", x"f7f1", 
            x"fb6c", x"fe27", x"00ad", x"03f1", 
            x"0703", x"0797", x"054f", x"027b", 
            x"0117", x"0100", x"01a6", x"036d", 
            x"0647", x"0889", x"08f1", x"0892", 
            x"08b0", x"084c", x"0609", x"02ca", 
            x"ffdd", x"fcf3", x"fa51", x"fa15", 
            x"fcc9", x"fee7", x"fcc0", x"f75a", 
            x"f326", x"f35f", x"f7d0", x"fd94", 
            x"0140", x"0198", x"006e", x"0079", 
            x"029a", x"04a7", x"0330", x"fdb0", 
            x"f7b1", x"f533", x"f708", x"fb4c", 
            x"0046", x"04e0", x"07df", x"0872", 
            x"077f", x"06b5", x"05af", x"02a6", 
            x"fde7", x"fa41", x"f9d4", x"fc5a", 
            x"0059", x"042a", x"0668", x"069d", 
            x"05ba", x"0501", x"0504", x"05c6", 
            x"0737", x"08a9", x"0877", x"0586", 
            x"01b7", x"00fa", x"0460", x"07f9", 
            x"0780", x"03e9", x"0191", x"0264", 
            x"0498", x"0670", x"07f7", x"08f8", 
            x"084c", x"05c0", x"02d8", x"01cb", 
            x"03c6", x"080f", x"0c33", x"0d88", 
            x"0b7c", x"07bb", x"0430", x"0247", 
            x"029c", x"045c", x"05bb", x"05a5", 
            x"04d7", x"04d0", x"057b", x"05a0", 
            x"0533", x"0549", x"060e", x"0619", 
            x"043e", x"011f", x"ff20", x"0019", 
            x"034a", x"0686", x"0896", x"0981", 
            x"093a", x"07bb", x"0661", x"0662", 
            x"0684", x"04ea", x"01ce", x"ff22", 
            x"fe15", x"fdf5", x"fddc", x"fe68", 
            x"004c", x"0341", x"06ca", x"0a22", 
            x"0bda", x"0ae8", x"0840", x"05a2", 
            x"032a", x"ffe4", x"fc3a", x"fa09", 
            x"f9ec", x"fa89", x"fb4b", x"fe16", 
            x"042f", x"0b11", x"0e70", x"0d06", 
            x"091a", x"0583", x"0352", x"0209", 
            x"0081", x"fe1a", x"fb6c", x"f983", 
            x"f8bc", x"f863", x"f7b1", x"f711", 
            x"f7a6", x"f94e", x"fa1d", x"f91a", 
            x"f82f", x"f94e", x"fae9", x"f9ec", 
            x"f666", x"f378", x"f2e8", x"f377", 
            x"f41a", x"f56e", x"f822", x"fbc0", 
            x"ff87", x"032d", x"0632", x"0778", 
            x"0664", x"0386", x"006b", x"fefd", 
            x"0059", x"038f", x"06ad", x"08e6", 
            x"0a39", x"09fa", x"0805", x"064c", 
            x"06d3", x"0836", x"0722", x"02b5", 
            x"fd44", x"f9b3", x"f979", x"fc3d", 
            x"0057", x"0454", x"07d5", x"0ad4", 
            x"0c3f", x"0a8c", x"0661", x"02a7", 
            x"00f9", x"00ec", x"020c", x"03c0", 
            x"0414", x"0186", x"fdcc", x"fca3", 
            x"ff51", x"02e6", x"0387", x"006b", 
            x"fcd1", x"fd04", x"0204", x"07f5", 
            x"0a15", x"0779", x"02fe", x"ff83", 
            x"fd92", x"fc95", x"fbca", x"faa0", 
            x"f905", x"f7fa", x"f89e", x"fa6c", 
            x"fb04", x"f92b", x"f761", x"f8ce", 
            x"fcaf", x"fee0", x"fd0e", x"f8e5", 
            x"f58b", x"f4fd", x"f7ea", x"fd67", 
            x"01de", x"013a", x"fc4a", x"f8e9", 
            x"fb0f", x"0024", x"02a2", x"0076", 
            x"fc32", x"f9c9", x"fb19", x"febb", 
            x"0134", x"0047", x"fd36", x"fa76", 
            x"f86d", x"f664", x"f50a", x"f52f", 
            x"f67c", x"f7c6", x"f7f4", x"f70a", 
            x"f6ab", x"f896", x"fbab", x"fc79", 
            x"f9ef", x"f6ac", x"f4db", x"f411", 
            x"f332", x"f244", x"f1e1", x"f250", 
            x"f37d", x"f4cc", x"f528", x"f42e", 
            x"f290", x"f0b0", x"ef19", x"ef51", 
            x"f266", x"f761", x"fb6a", x"fbe5", 
            x"f935", x"f5b3", x"f363", x"f322", 
            x"f46f", x"f58f", x"f4f2", x"f365", 
            x"f34d", x"f5b7", x"f909", x"fb58", 
            x"fc7e", x"fd58", x"fe3c", x"fee0", 
            x"ff60", x"0087", x"0240", x"032c", 
            x"02ab", x"026f", x"044d", x"0700", 
            x"07b4", x"05c6", x"02ae", x"ffe8", 
            x"fdff", x"fce1", x"fca0", x"fd89", 
            x"ff86", x"01ff", x"0443", x"05e2", 
            x"0725", x"084d", x"089c", x"06ce", 
            x"02e2", x"fefc", x"fd92", x"ff76", 
            x"03b3", x"08db", x"0db0", x"10f3", 
            x"114a", x"0e2c", x"0934", x"0531", 
            x"044a", x"06e2", x"0aeb", x"0d7a", 
            x"0e11", x"0f2a", x"12c2", x"16cf", 
            x"1739", x"131c", x"0d54", x"088e", 
            x"0578", x"0431", x"049c", x"05c0", 
            x"067f", x"0656", x"0529", x"0359", 
            x"0279", x"03fa", x"0678", x"075f", 
            x"069c", x"05b1", x"0519", x"04a4", 
            x"04c9", x"0673", x"092c", x"0ab9", 
            x"09ee", x"08e9", x"0a8b", x"0f05", 
            x"1385", x"1507", x"133d", x"1034", 
            x"0db3", x"0c4e", x"0c74", x"0e0a", 
            x"0f28", x"0d7a", x"0996", x"0613", 
            x"0430", x"035a", x"02b7", x"01ce", 
            x"0068", x"fed7", x"fe22", x"ff28", 
            x"018c", x"0407", x"055a", x"04f4", 
            x"0394", x"0284", x"01b7", x"0083", 
            x"0000", x"0308", x"0a5d", x"1240", 
            x"15fc", x"146a", x"0ff7", x"0b7c", 
            x"0814", x"05ae", x"048e", x"0553", 
            x"07ae", x"0a05", x"0a36", x"06ce", 
            x"009c", x"fa3e", x"f621", x"f4c8", 
            x"f514", x"f632", x"f856", x"fbc2", 
            x"ffe8", x"0374", x"0460", x"014b", 
            x"fb10", x"f48d", x"efdc", x"ecb4", 
            x"ea4a", x"e8fd", x"e91e", x"e9ee", 
            x"eaf7", x"ec7e", x"ee8b", x"f033", 
            x"f122", x"f244", x"f3c5", x"f486", 
            x"f3db", x"f26b", x"f11f", x"f097", 
            x"f13e", x"f328", x"f58d", x"f719", 
            x"f83b", x"fbd7", x"0322", x"0a2f", 
            x"0ba1", x"0772", x"0314", x"0224", 
            x"0254", x"0030", x"fd0c", x"fcf4", 
            x"00ea", x"056c", x"0685", x"03f7", 
            x"00a3", x"ff78", x"0084", x"0131", 
            x"ffc0", x"fcf9", x"fa4e", x"f7fe", 
            x"f5e1", x"f459", x"f3fc", x"f488", 
            x"f507", x"f4fb", x"f4eb", x"f54b", 
            x"f5b1", x"f618", x"f727", x"f946", 
            x"fb98", x"fc84", x"fbad", x"fac0", 
            x"fb7b", x"fdb5", x"ffe5", x"00fc", 
            x"011b", x"009b", x"ffeb", x"ffe6", 
            x"016e", x"040a", x"069a", x"08eb", 
            x"0aab", x"0a7d", x"07c6", x"04c7", 
            x"042c", x"0578", x"0639", x"05e3", 
            x"05e8", x"06b3", x"0706", x"0617", 
            x"0433", x"0197", x"fead", x"fcbb", 
            x"fc30", x"fb49", x"f927", x"f841", 
            x"fb0e", x"ffd0", x"01fe", x"ffcc", 
            x"fbe7", x"f98d", x"f8d4", x"f802", 
            x"f6d3", x"f6a4", x"f881", x"fc08", 
            x"ff95", x"00ee", x"ff0a", x"fb78", 
            x"f8f6", x"f80d", x"f6cf", x"f471", 
            x"f335", x"f498", x"f6b7", x"f792", 
            x"f7ed", x"f909", x"fa2e", x"fa87", 
            x"faaf", x"fac2", x"fa2a", x"f9a6", 
            x"fa4a", x"fba5", x"fc9f", x"fdb7", 
            x"003b", x"039f", x"0581", x"0441", 
            x"005f", x"fb99", x"f7d6", x"f66d", 
            x"f7be", x"fac7", x"fdd9", x"ffa1", 
            x"0011", x"00b3", x"0305", x"0654", 
            x"083d", x"0793", x"053e", x"026f", 
            x"ffe3", x"fe98", x"ff29", x"0165"
        ),
        -- Block 20
        (
            x"054d", x"0a84", x"0ecf", x"0fdb", 
            x"0e2d", x"0cb6", x"0d55", x"0ee6", 
            x"0f7d", x"0ed6", x"0e2b", x"0dca", 
            x"0c94", x"09f8", x"075b", x"06a3", 
            x"0770", x"06a8", x"0270", x"fd72", 
            x"fb69", x"fc49", x"fd10", x"fc44", 
            x"fad6", x"f9eb", x"f92b", x"f6a5", 
            x"f106", x"eaa3", x"e82e", x"eb3d", 
            x"f014", x"f1e6", x"f06d", x"efd1", 
            x"f2a5", x"f737", x"fac4", x"fce5", 
            x"fed6", x"00e5", x"0243", x"02bd", 
            x"03b7", x"0664", x"09df", x"0cb5", 
            x"0efa", x"10c4", x"108e", x"0da9", 
            x"0a5c", x"097a", x"0a83", x"0aee", 
            x"09cb", x"0812", x"06bb", x"0624", 
            x"063b", x"0637", x"0524", x"02d3", 
            x"0049", x"ff2d", x"0067", x"0378", 
            x"06ec", x"099e", x"0b68", x"0cce", 
            x"0e60", x"1011", x"10ba", x"0e95", 
            x"0915", x"02ad", x"ff13", x"ff47", 
            x"0149", x"0370", x"053d", x"05b5", 
            x"0446", x"02fc", x"046c", x"07c9", 
            x"0944", x"0628", x"ffaf", x"f9f5", 
            x"f84f", x"fad4", x"ff49", x"02d7", 
            x"036c", x"011c", x"fde6", x"fc7d", 
            x"fe3e", x"01cd", x"049e", x"058d", 
            x"04f1", x"0360", x"0208", x"0248", 
            x"0434", x"06b2", x"08c8", x"0a14", 
            x"0a31", x"0904", x"0739", x"05cd", 
            x"0523", x"058d", x"077e", x"09ef", 
            x"0a13", x"0612", x"0004", x"fc98", 
            x"fdd4", x"00ce", x"00fb", x"fd6a", 
            x"f9ff", x"faf5", x"fff7", x"052d", 
            x"07bf", x"0752", x"04c7", x"01c5", 
            x"0087", x"023e", x"053b", x"0695", 
            x"05d2", x"04f9", x"0551", x"05ef", 
            x"0625", x"06de", x"08a1", x"09aa", 
            x"0775", x"0238", x"fd3c", x"fb05", 
            x"fb63", x"fd1e", x"ff4a", x"0039", 
            x"fde8", x"f8f9", x"f4fe", x"f4e2", 
            x"f82f", x"fc86", x"0000", x"0195", 
            x"00fb", x"ff2d", x"fd5b", x"fbcd", 
            x"fa97", x"fa08", x"f976", x"f7b6", 
            x"f598", x"f5f3", x"f9b5", x"fe29", 
            x"007b", x"0065", x"ff3c", x"fe41", 
            x"fd89", x"fbd6", x"f83f", x"f3c3", 
            x"f0ff", x"f194", x"f3e3", x"f54e", 
            x"f592", x"f634", x"f761", x"f75b", 
            x"f502", x"f162", x"eecd", x"eede", 
            x"f0ce", x"f1aa", x"efdd", x"ed97", 
            x"ee8c", x"f381", x"f96b", x"fd17", 
            x"fe5c", x"ffb7", x"033b", x"0856", 
            x"0c2c", x"0c60", x"0995", x"0656", 
            x"03a5", x"00b9", x"fd52", x"fa6e", 
            x"f99c", x"fb68", x"fedc", x"0205", 
            x"0353", x"0276", x"0030", x"fd5b", 
            x"fa56", x"f673", x"f1c6", x"ef12", 
            x"f0e4", x"f4f2", x"f61a", x"f39a", 
            x"f268", x"f61a", x"fbcb", x"fe67", 
            x"fdc2", x"fd37", x"fd46", x"fc41", 
            x"fb2c", x"fd69", x"0368", x"0940", 
            x"0b91", x"0ae3", x"0931", x"06ae", 
            x"027e", x"fcff", x"f8a3", x"f814", 
            x"fad4", x"fd61", x"fd9c", x"fd36", 
            x"fe20", x"ff20", x"fda5", x"f995", 
            x"f58d", x"f357", x"f28a", x"f2c8", 
            x"f537", x"fa73", x"0078", x"0406", 
            x"038d", x"009d", x"fecf", x"00b2", 
            x"0564", x"0903", x"084c", x"03f3", 
            x"0007", x"ff99", x"01cd", x"03ae", 
            x"036d", x"0205", x"0298", x"073f", 
            x"0db1", x"10b5", x"0e28", x"094d", 
            x"062c", x"051c", x"0437", x"02cb", 
            x"01a9", x"01cf", x"0383", x"05fc", 
            x"06e6", x"045b", x"0083", x"002f", 
            x"0445", x"0858", x"0911", x"082c", 
            x"088c", x"0a16", x"0af3", x"09f2", 
            x"06b7", x"01b6", x"fcc9", x"f9da", 
            x"f989", x"fb0b", x"fd96", x"00a5", 
            x"0363", x"0520", x"0640", x"0788", 
            x"088f", x"07f5", x"054a", x"01c6", 
            x"ff04", x"fe84", x"00bd", x"0431", 
            x"0655", x"05d7", x"037a", x"00b3", 
            x"fddd", x"faba", x"f868", x"f830", 
            x"f8f7", x"f7f0", x"f461", x"f107", 
            x"f104", x"f3a5", x"f52d", x"f430", 
            x"f331", x"f41a", x"f66c", x"f95b", 
            x"fc1e", x"fd29", x"fc4f", x"fbeb", 
            x"fd2e", x"fe5b", x"fe0f", x"fd40", 
            x"fcec", x"fc4e", x"fa6d", x"f7f4", 
            x"f652", x"f664", x"f817", x"fa64", 
            x"fc07", x"fce5", x"fe26", x"00b2", 
            x"03da", x"0664", x"07b7", x"06ac", 
            x"0220", x"fbc8", x"f7e6", x"f84b", 
            x"fae9", x"fd45", x"feff", x"00dd", 
            x"0359", x"0630", x"07bb", x"0628", 
            x"01e0", x"fd61", x"fae4", x"fb61", 
            x"fea1", x"02d3", x"057e", x"05c9", 
            x"04f4", x"03bb", x"0142", x"fda3", 
            x"faee", x"fa56", x"fab7", x"fbe1", 
            x"ff7b", x"0514", x"08e2", x"0829", 
            x"04ae", x"0239", x"02c9", x"04bc", 
            x"048f", x"015e", x"fe62", x"fe80", 
            x"0075", x"0144", x"0082", x"ffe1", 
            x"0015", x"0021", x"ff54", x"fe2a", 
            x"fd5b", x"fd30", x"fd8f", x"fe3d", 
            x"ffb4", x"0270", x"053d", x"0694", 
            x"0729", x"08b7", x"0aa1", x"0a6f", 
            x"0726", x"039f", x"0402", x"089d", 
            x"0d69", x"0eb3", x"0c27", x"0825", 
            x"05fb", x"06dd", x"0886", x"07f5", 
            x"0518", x"0222", x"00cc", x"0127", 
            x"026a", x"0332", x"018b", x"fd4f", 
            x"f956", x"f88e", x"fa53", x"fb3f", 
            x"f9fd", x"f8ad", x"f8ca", x"f911", 
            x"f877", x"f7eb", x"f7cc", x"f700", 
            x"f57c", x"f4f2", x"f646", x"f83f", 
            x"f987", x"fa11", x"fa40", x"f9eb", 
            x"f953", x"f9f4", x"fdc7", x"048f", 
            x"0b20", x"0e99", x"0f20", x"0e65", 
            x"0d11", x"0aa2", x"06c5", x"0257", 
            x"ff45", x"ffcf", x"0499", x"0adb", 
            x"0e42", x"0de3", x"0d0c", x"0ea7", 
            x"1170", x"1222", x"0fc0", x"0bc8", 
            x"08c9", x"0890", x"09f5", x"09a4", 
            x"0642", x"01b7", x"fe04", x"fb52", 
            x"f974", x"f8ce", x"f91d", x"f986", 
            x"fa22", x"fb77", x"fcac", x"fce2", 
            x"fcd0", x"fd59", x"fe56", x"ffa8", 
            x"0178", x"02dc", x"0297", x"0175", 
            x"0172", x"02b4", x"045a", x"06bf", 
            x"0a01", x"0c1d", x"0bc0", x"0ab1", 
            x"0b88", x"0e7b", x"1152", x"11af", 
            x"0e48", x"07d4", x"0176", x"fe6e", 
            x"fec1", x"ffeb", x"007d", x"0115", 
            x"0281", x"040a", x"034b", x"ff17", 
            x"f9e3", x"f721", x"f6ea", x"f604", 
            x"f2d9", x"f072", x"f22f", x"f718", 
            x"fb46", x"fce4", x"fd6d", x"fe97", 
            x"ffd1", x"0006", x"fff5", x"015c", 
            x"0415", x"0564", x"03a2", x"008b", 
            x"fe8c", x"fe00", x"fea9", x"00ee", 
            x"0483", x"072b", x"06cc", x"04a4", 
            x"040d", x"067d", x"09ee", x"0ab3", 
            x"06f2", x"00fe", x"fd79", x"fdd6", 
            x"fe05", x"fa85", x"f5b8", x"f39e", 
            x"f46a", x"f5bf", x"f634", x"f5c4", 
            x"f4f6", x"f4df", x"f673", x"f847", 
            x"f752", x"f32e", x"ef17", x"ee36", 
            x"f084", x"f3d1", x"f62d", x"f69e", 
            x"f591", x"f4b3", x"f54d", x"f6da", 
            x"f7ac", x"f705", x"f64b", x"f793", 
            x"fb46", x"ffde", x"03b3", x"05cd", 
            x"05be", x"0402", x"0292", x"0375", 
            x"0663", x"084e", x"071e", x"0512", 
            x"0582", x"07c7", x"08a4", x"06f4", 
            x"03e5", x"0084", x"fd9f", x"fcd6", 
            x"ff46", x"0322", x"049b", x"01eb", 
            x"fd7b", x"fb13", x"fb66", x"fb6b", 
            x"f8fd", x"f61c", x"f546", x"f57a", 
            x"f501", x"f4cd", x"f610", x"f77d", 
            x"f6c5", x"f30b", x"edc3", x"ea3f", 
            x"eb47", x"f02e", x"f633", x"fbec", 
            x"0126", x"048e", x"04a2", x"0296", 
            x"00de", x"ff51", x"fbc1", x"f68c", 
            x"f2f9", x"f34b", x"f655", x"f917", 
            x"f9ea", x"f90f", x"f836", x"f987", 
            x"fd84", x"01a1", x"032f", x"025b", 
            x"011a", x"0095", x"00bb", x"0086", 
            x"fe71", x"fa68", x"f66a", x"f4d1", 
            x"f6c4", x"fb91", x"006c", x"0240", 
            x"0053", x"fd12", x"fb8c", x"fc8d", 
            x"fe5f", x"feef", x"fde2", x"fca4", 
            x"fca3", x"fe0a", x"0058", x"02ef", 
            x"0507", x"05e0", x"04a9", x"00d6", 
            x"fbef", x"f923", x"f9bb", x"fc20", 
            x"fe62", x"005c", x"030e", x"0685", 
            x"08dc", x"08ec", x"086a", x"09d7", 
            x"0d80", x"1131", x"12f1", x"1389", 
            x"1553", x"1827", x"1880", x"1425", 
            x"0d9a", x"0980", x"09b6", x"0c30", 
            x"0e31", x"0f18", x"0fbc", x"1080", 
            x"111a", x"113f", x"107d", x"0e35", 
            x"0ad3", x"0874", x"08f5", x"0b3e", 
            x"0bd7", x"08fd", x"0430", x"fff5", 
            x"fdbe", x"fd89", x"fda8", x"fc4b", 
            x"fa78", x"fb74", x"005f", x"06a6", 
            x"0abc", x"0b11", x"0845", x"03e9", 
            x"0014", x"fe7a", x"feab", x"fe47", 
            x"fc75", x"fb4b", x"fc20", x"fd5d", 
            x"fd3e", x"fba2", x"f9f3", x"fa27", 
            x"fcca", x"0048", x"036c", x"06aa", 
            x"0a29", x"0bfd", x"0a52", x"05ff", 
            x"01fb", x"007f", x"017d", x"0312", 
            x"0366", x"0237", x"0106", x"0159", 
            x"02d0", x"045d", x"065f", x"08fd", 
            x"0a65", x"094d", x"071f", x"0622", 
            x"060c", x"041e", x"feb4", x"f814", 
            x"f45a", x"f51b", x"f82d", x"fa00", 
            x"f93e", x"f7a1", x"f6fa", x"f71b", 
            x"f772", x"f7dd", x"f7ca", x"f6e2", 
            x"f637", x"f775", x"fafc", x"ff80", 
            x"03b5", x"0758", x"09b3", x"09d1", 
            x"0812", x"061d", x"052f", x"0539", 
            x"054a", x"0526", x"05f1", x"08b4", 
            x"0cfa", x"11c7", x"1626", x"1857", 
            x"174f", x"146c", x"1155", x"0dd8", 
            x"094d", x"0499", x"014d", x"ff28", 
            x"fccb", x"fae5", x"fb3f", x"fd41", 
            x"fde4", x"fb5d", x"f6eb", x"f308", 
            x"f0d0", x"f03b", x"f0c8", x"f162", 
            x"f256", x"f578", x"fa39", x"fcf3", 
            x"fbee", x"fa0e", x"fb02", x"fde8", 
            x"ff0d", x"fdf9", x"fe12", x"01a8", 
            x"076a", x"0c02", x"0cef", x"0a66", 
            x"077f", x"06f0", x"0764", x"05ad", 
            x"0278", x"01b1", x"0405", x"05ad", 
            x"0465", x"01a6", x"fea7", x"fb33", 
            x"f84d", x"f7dd", x"f956", x"f995", 
            x"f6d3", x"f2c2", x"f055", x"f15c", 
            x"f58d", x"fa93", x"fdd3", x"fe9e", 
            x"fdf9", x"fcce", x"faa0", x"f677", 
            x"f182", x"ef2f", x"f184", x"f68a", 
            x"fa29", x"fae9", x"fb3d", x"fd0b", 
            x"ff48", x"00eb", x"0251", x"02dc", 
            x"00e2", x"fd30", x"fb6c", x"fdad", 
            x"01a1", x"039b", x"02be", x"018e", 
            x"02ef", x"0743", x"0b9c", x"0c51", 
            x"08b1", x"03b7", x"0112", x"01fe", 
            x"047d", x"050a", x"022a", x"fe44", 
            x"fc1a", x"faea", x"f934", x"f823", 
            x"f8fc", x"fa27", x"f98a", x"f80c", 
            x"f86b", x"fab3", x"fc1c", x"fb01", 
            x"f836", x"f56d", x"f433", x"f532", 
            x"f76e", x"f95e", x"fb6b", x"ff30", 
            x"03d5", x"0619", x"04bb", x"01ca", 
            x"ffa5", x"feb2", x"fdcb", x"fbb0", 
            x"f87d", x"f60b", x"f6a2", x"faa9", 
            x"ffc2", x"032e", x"0528", x"076e", 
            x"0980", x"0937", x"06ee", x"0558", 
            x"04df", x"02f8", x"fe62", x"f944", 
            x"f6a5", x"f720", x"f8cd", x"f9cb", 
            x"f9e3", x"f917", x"f6d1", x"f34f", 
            x"f078", x"efe9", x"f0f4", x"f1aa", 
            x"f13d", x"f0b4", x"f1e2", x"f571", 
            x"f9f6", x"fd46", x"feb0", x"ff3d", 
            x"ffdc", x"004d", x"0027", x"001a", 
            x"0164", x"03aa", x"0490", x"0278", 
            x"ff4a", x"fdde", x"fecb", x"0130", 
            x"041c", x"05f7", x"0517", x"01d8", 
            x"fec4", x"fdb2", x"fdd7", x"fd8f", 
            x"fc43", x"fa4d", x"f863", x"f775", 
            x"f796", x"f78b", x"f61a", x"f350", 
            x"f085", x"efa7", x"f1b8", x"f555", 
            x"f7ff", x"f803", x"f5f2", x"f46a", 
            x"f510", x"f6a8", x"f7e3", x"f945"
        ),
        -- Block 19
        (
            x"faa4", x"fa2b", x"f793", x"f5c6", 
            x"f6ab", x"f8ea", x"faec", x"fd65", 
            x"0108", x"04d0", x"0775", x"0904", 
            x"0aa1", x"0cf3", x"0f58", x"10c5", 
            x"10af", x"0f6b", x"0e16", x"0dbe", 
            x"0ddf", x"0c85", x"0903", x"04e4", 
            x"01e9", x"006e", x"0004", x"0078", 
            x"01be", x"02e7", x"01fe", x"fe1e", 
            x"f983", x"f7d6", x"fa21", x"fd64", 
            x"fe84", x"fe09", x"fe88", x"00df", 
            x"0383", x"04a9", x"0412", x"02cd", 
            x"01f4", x"022b", x"035b", x"04e6", 
            x"0617", x"06a1", x"077d", x"0a23", 
            x"0e4d", x"1199", x"122a", x"109a", 
            x"0efa", x"0e4c", x"0dba", x"0c31", 
            x"09fd", x"089d", x"096c", x"0c21", 
            x"0ef1", x"1029", x"0f7d", x"0d56", 
            x"0a66", x"07c9", x"060d", x"0453", 
            x"024d", x"0161", x"023b", x"035b", 
            x"0327", x"02b2", x"0408", x"06a3", 
            x"0769", x"050b", x"0291", x"03ae", 
            x"083c", x"0c91", x"0cdc", x"0866", 
            x"02dd", x"007b", x"01b7", x"040d", 
            x"050a", x"03fa", x"0236", x"0231", 
            x"0529", x"09bb", x"0d82", x"0f90", 
            x"106f", x"101e", x"0dbe", x"09aa", 
            x"05e1", x"03e2", x"0386", x"0399", 
            x"030a", x"0181", x"ffbb", x"fec7", 
            x"ff17", x"0062", x"0285", x"05e8", 
            x"09c3", x"0b91", x"09bc", x"055d", 
            x"00f3", x"fe72", x"fea6", x"00e8", 
            x"039f", x"05a8", x"0624", x"03ff", 
            x"ffc7", x"fca8", x"fdc5", x"025c", 
            x"05ed", x"051b", x"0179", x"ff26", 
            x"ff46", x"fe66", x"f963", x"f243", 
            x"ee0f", x"ef54", x"f45c", x"f916", 
            x"fa7b", x"f8b0", x"f663", x"f677", 
            x"f975", x"fc7d", x"fc42", x"f90f", 
            x"f6c2", x"f7dd", x"fa50", x"faee", 
            x"f945", x"f689", x"f31e", x"eff0", 
            x"ef35", x"f17f", x"f443", x"f4e8", 
            x"f3ac", x"f2c4", x"f350", x"f406", 
            x"f2ca", x"f01a", x"efb4", x"f3dd", 
            x"f903", x"f9cb", x"f61c", x"f32a", 
            x"f589", x"fc40", x"020a", x"036a", 
            x"023e", x"0276", x"054b", x"08c6", 
            x"0a88", x"0996", x"0642", x"018c", 
            x"fd08", x"fa5c", x"fa12", x"fb89", 
            x"fdbd", x"ff7a", x"fef1", x"fa8d", 
            x"f47e", x"f1e5", x"f450", x"f779", 
            x"f7ff", x"f796", x"f88c", x"fa17", 
            x"fb12", x"fcfa", x"00b4", x"02e7", 
            x"ffff", x"fa4c", x"f7a1", x"f9b7", 
            x"fd2c", x"ff44", x"0067", x"014d", 
            x"0158", x"009e", x"00e1", x"02d7", 
            x"04ef", x"067f", x"0930", x"0d47", 
            x"0f93", x"0d09", x"06f9", x"01a2", 
            x"ffb6", x"000b", x"ff79", x"fc48", 
            x"f809", x"f5b9", x"f68b", x"f95f", 
            x"fc41", x"fda4", x"fd23", x"fbce", 
            x"fb92", x"fd44", x"0041", x"0433", 
            x"0935", x"0d1d", x"0c13", x"0604", 
            x"0016", x"fee6", x"020c", x"05b9", 
            x"063d", x"029e", x"fcb9", x"f74d", 
            x"f421", x"f35c", x"f42a", x"f632", 
            x"fa38", x"000f", x"0474", x"03a0", 
            x"fe43", x"f89d", x"f4cb", x"f1b4", 
            x"ee81", x"ec98", x"ee0f", x"f2eb", 
            x"f9b8", x"0118", x"06cc", x"088b", 
            x"0719", x"055c", x"03d4", x"00d2", 
            x"fe09", x"ffea", x"0645", x"0b89", 
            x"0cbb", x"0ca2", x"0e44", x"1066", 
            x"0fda", x"0c18", x"07f5", x"0618", 
            x"06a3", x"0802", x"08b7", x"0869", 
            x"07fe", x"083c", x"08bb", x"0917", 
            x"09c1", x"0a53", x"093f", x"0751", 
            x"0722", x"085e", x"07e7", x"04fc", 
            x"0266", x"0221", x"0354", x"03e7", 
            x"029d", x"0027", x"fe5c", x"fe18", 
            x"fe4c", x"fcee", x"f910", x"f46b", 
            x"f190", x"f0b9", x"f07b", x"f091", 
            x"f229", x"f5d4", x"f9c9", x"fa77", 
            x"f6af", x"f228", x"f18f", x"f551", 
            x"f9d5", x"fbe4", x"fbb0", x"fc5c", 
            x"00a6", x"0750", x"0bb4", x"0a53", 
            x"0535", x"02ab", x"0670", x"0d9f", 
            x"129a", x"128e", x"0e7a", x"09a6", 
            x"07bc", x"092e", x"0a33", x"0791", 
            x"02db", x"00f4", x"040c", x"083b", 
            x"086c", x"054b", x"0360", x"0392", 
            x"0241", x"fd77", x"f7f1", x"f504", 
            x"f456", x"f391", x"f1d9", x"efc2", 
            x"ee3b", x"ee42", x"efc7", x"f127", 
            x"f1be", x"f365", x"f776", x"fd31", 
            x"036d", x"08d1", x"0aaa", x"07b7", 
            x"03c2", x"036d", x"054d", x"04e1", 
            x"0292", x"02e4", x"0687", x"0944", 
            x"08c9", x"0730", x"0612", x"0406", 
            x"0071", x"fd71", x"fd11", x"ff74", 
            x"02f3", x"0508", x"03da", x"005e", 
            x"fd5c", x"fb83", x"f85e", x"f274", 
            x"ebf5", x"e868", x"e960", x"ed8f", 
            x"f2d6", x"f830", x"fcf6", x"0023", 
            x"00ef", x"ffd1", x"fe84", x"fe85", 
            x"ffba", x"009a", x"0052", x"0001", 
            x"0176", x"045e", x"06cd", x"0841", 
            x"09de", x"0b84", x"0b98", x"0a36", 
            x"0a37", x"0d2c", x"10c1", x"11ae", 
            x"0fc1", x"0d8d", x"0d3a", x"0dfa", 
            x"0d6b", x"0bb0", x"0b4e", x"0ccd", 
            x"0d6f", x"0b99", x"09d4", x"0a7d", 
            x"0b0f", x"0785", x"007f", x"fa90", 
            x"f8ec", x"faaf", x"fca7", x"fc01", 
            x"f83b", x"f3f7", x"f262", x"f323", 
            x"f350", x"f246", x"f28a", x"f619", 
            x"fc2e", x"02f1", x"0899", x"0b82", 
            x"0b06", x"07d6", x"0366", x"ff5a", 
            x"fd36", x"fd60", x"fe61", x"ff2c", 
            x"014c", x"05e3", x"0a42", x"0acc", 
            x"0886", x"07a0", x"08e7", x"08fd", 
            x"0614", x"027b", x"015e", x"028f", 
            x"035c", x"0285", x"0150", x"0164", 
            x"02c8", x"03db", x"0353", x"0235", 
            x"0225", x"02d9", x"037e", x"04cc", 
            x"0701", x"07e4", x"0577", x"0127", 
            x"fe2e", x"fd6f", x"fcfd", x"fb04", 
            x"f818", x"f6cf", x"f981", x"ff25", 
            x"0320", x"0237", x"fe2c", x"fac3", 
            x"f97b", x"f95a", x"f92c", x"f8d6", 
            x"f932", x"fac2", x"fc6d", x"fc7d", 
            x"fb68", x"fb49", x"fc04", x"fb9d", 
            x"fa54", x"fac3", x"fdcb", x"013f", 
            x"02e7", x"02d9", x"02ee", x"04c3", 
            x"080b", x"0a3b", x"091e", x"0653", 
            x"0591", x"0651", x"03ad", x"fbeb", 
            x"f45f", x"f326", x"f7b9", x"fcc1", 
            x"feb4", x"fe6a", x"fe6f", x"ff95", 
            x"0004", x"fe2c", x"fae7", x"f869", 
            x"f827", x"f9ad", x"fafe", x"fb2e", 
            x"fb94", x"fc89", x"fbfe", x"f93d", 
            x"f662", x"f523", x"f4ff", x"f5aa", 
            x"f7ee", x"fb5a", x"fe4e", x"0087", 
            x"0374", x"0661", x"04fb", x"fd77", 
            x"f5a6", x"f4bb", x"fad2", x"02a4", 
            x"0895", x"0c51", x"0e00", x"0d16", 
            x"0965", x"0413", x"fede", x"fb05", 
            x"f89c", x"f72f", x"f7c1", x"fc1b", 
            x"0261", x"0513", x"024d", x"fecf", 
            x"fe49", x"fdd8", x"f972", x"f302", 
            x"f064", x"f3d9", x"f9a9", x"fccd", 
            x"fc99", x"fc59", x"fe42", x"0125", 
            x"0324", x"0473", x"062d", x"080f", 
            x"093b", x"09d5", x"0a4c", x"09e9", 
            x"07e8", x"04f1", x"01ae", x"fe50", 
            x"fb52", x"f97f", x"f9ab", x"fbf4", 
            x"fefb", x"00cf", x"0117", x"0184", 
            x"034d", x"0584", x"06ca", x"06be", 
            x"0538", x"026b", x"0021", x"00a5", 
            x"030d", x"0303", x"fe3b", x"f791", 
            x"f2ce", x"f11c", x"f2da", x"f7f4", 
            x"fe16", x"01ee", x"029f", x"01f1", 
            x"0207", x"0380", x"0501", x"0461", 
            x"00e9", x"fcf7", x"fb77", x"fc03", 
            x"fbd9", x"fa89", x"fa35", x"fbb3", 
            x"fdd6", x"ffe1", x"0214", x"0423", 
            x"04b5", x"03be", x"035f", x"04b1", 
            x"059a", x"03f0", x"0167", x"0172", 
            x"03f9", x"0548", x"034b", x"00a6", 
            x"010b", x"03b8", x"0505", x"0470", 
            x"04da", x"07cb", x"0b34", x"0bda", 
            x"08fe", x"04f4", x"0273", x"01c7", 
            x"0112", x"febd", x"fb1e", x"f794", 
            x"f474", x"f155", x"ef11", x"efc8", 
            x"f404", x"f9a4", x"fe38", x"00c6", 
            x"01c4", x"0234", x"0210", x"ffc7", 
            x"fb4f", x"f7a8", x"f74f", x"f9ea", 
            x"fded", x"0229", x"058c", x"06fd", 
            x"0686", x"058c", x"04a0", x"02c8", 
            x"0054", x"ffc1", x"025b", x"06a5", 
            x"0b26", x"0fcb", x"13fe", x"15dc", 
            x"13c0", x"0d76", x"04b3", x"fcd8", 
            x"f8d1", x"f8ca", x"f9f7", x"f9e4", 
            x"f916", x"f928", x"fa69", x"fc2a", 
            x"fdd6", x"fe41", x"fc43", x"f96d", 
            x"f8f8", x"fb67", x"fe90", x"0191", 
            x"0555", x"09a4", x"0be2", x"0a5b", 
            x"068c", x"02e8", x"0004", x"fd91", 
            x"fc3f", x"fd15", x"ffbd", x"0298", 
            x"0439", x"046c", x"042a", x"03fe", 
            x"0336", x"0129", x"fea5", x"fdb7", 
            x"ff77", x"0240", x"03bf", x"03c1", 
            x"0383", x"0396", x"03c7", x"0457", 
            x"05a3", x"075a", x"0849", x"073d", 
            x"0445", x"0101", x"fedd", x"fe68", 
            x"0041", x"03c1", x"06c6", x"08b7", 
            x"0a96", x"0b95", x"0a1b", x"0858", 
            x"0a44", x"0e0f", x"0c9a", x"0405", 
            x"fbad", x"fa15", x"fbff", x"faa6", 
            x"f664", x"f442", x"f49b", x"f42e", 
            x"f3cb", x"f6d2", x"fb84", x"fcb7", 
            x"fa43", x"f892", x"f941", x"f9f6", 
            x"f9a9", x"fa10", x"fb87", x"fbf5", 
            x"fafe", x"fae4", x"fbfb", x"fbd1", 
            x"fa1f", x"f9ef", x"fc91", x"ffbc", 
            x"0190", x"0213", x"0067", x"fb8f", 
            x"f611", x"f3c2", x"f3e5", x"f291", 
            x"ef92", x"ef37", x"f314", x"f6e0", 
            x"f66f", x"f35a", x"f1ce", x"f1f1", 
            x"f0f7", x"ee6f", x"ebdb", x"e98d", 
            x"e7d4", x"e89c", x"ecc3", x"f21b", 
            x"f616", x"f8c5", x"fc18", x"0107", 
            x"05cd", x"073f", x"0464", x"003f", 
            x"fe3f", x"fe14", x"fd2f", x"fb31", 
            x"fa66", x"fbc3", x"fdc2", x"ffb4", 
            x"027a", x"0480", x"02f4", x"ffb3", 
            x"ff35", x"0170", x"027d", x"009b", 
            x"fda9", x"fbd8", x"fbf3", x"fdc6", 
            x"ff94", x"ff53", x"fe10", x"fe7e", 
            x"ffb2", x"fdcd", x"f828", x"f337", 
            x"f38c", x"f870", x"fccf", x"fcd0", 
            x"f95e", x"f69e", x"f772", x"fab0", 
            x"fd4a", x"fec8", x"0161", x"0566", 
            x"07c7", x"0674", x"037f", x"0257", 
            x"03a7", x"051d", x"046e", x"0233", 
            x"0166", x"041c", x"0904", x"0c9a", 
            x"0cf5", x"0b98", x"0ac9", x"0a92", 
            x"0969", x"0631", x"01ba", x"fed8", 
            x"0005", x"0433", x"0745", x"069a", 
            x"0486", x"05ea", x"0b4a", x"0f56", 
            x"0eba", x"0c90", x"0b4f", x"0889", 
            x"031e", x"feae", x"fdf1", x"ff09", 
            x"ffb9", x"00e8", x"03e4", x"07e7", 
            x"0bb8", x"0e79", x"0f2c", x"0d5b", 
            x"09bf", x"05f4", x"02f3", x"00e1", 
            x"0089", x"026e", x"047b", x"043d", 
            x"02eb", x"0389", x"05ec", x"06c0", 
            x"048c", x"0195", x"0004", x"ff4d", 
            x"feb0", x"ff4b", x"01d2", x"0494", 
            x"0523", x"034f", x"0105", x"ff95", 
            x"fed0", x"febb", x"ff6d", x"ffe2", 
            x"fedf", x"fca8", x"fb41", x"fcee", 
            x"01f8", x"081b", x"0bc6", x"0a72", 
            x"05ae", x"0224", x"02c1", x"0685", 
            x"0ac6", x"0d9f", x"0eb8", x"0eaa", 
            x"0d95", x"0ab3", x"05cd", x"0113", 
            x"ff9d", x"00fd", x"00e3", x"fd19", 
            x"f8bf", x"f7e2", x"fa5d", x"fc80", 
            x"fb8b", x"f844", x"f54c", x"f38e", 
            x"f23c", x"f176", x"f30a", x"f853", 
            x"ff2a", x"0278", x"ffb2", x"fb1d", 
            x"fb0c", x"ff2f", x"0159", x"fe4d", 
            x"f949", x"f773", x"fa16", x"fd54", 
            x"fd6a", x"fc66", x"ff01", x"04bd", 
            x"07b6", x"04f3", x"0031", x"fe04", 
            x"fe78", x"fee6", x"fdd7", x"fbcd", 
            x"fa1d", x"f9be", x"fa9e", x"fbea"
        ),
        -- Block 18
        (
            x"fd38", x"ff57", x"030d", x"06a8", 
            x"0758", x"050e", x"02ea", x"03aa", 
            x"0717", x"0a58", x"0a6c", x"07bf", 
            x"0620", x"073f", x"07d6", x"04d7", 
            x"009b", x"ffbf", x"02c6", x"05b8", 
            x"0512", x"00c3", x"fb1b", x"f74a", 
            x"f7e1", x"fc37", x"008b", x"01fd", 
            x"0188", x"0194", x"01f7", x"00b9", 
            x"fdcb", x"fb86", x"fb19", x"fb02", 
            x"fa4c", x"faee", x"fe90", x"031e", 
            x"05bd", x"0700", x"0931", x"0bbc", 
            x"0b05", x"062e", x"0196", x"00a3", 
            x"00dc", x"fe74", x"fb00", x"fb00", 
            x"fe4f", x"003c", x"ff0e", x"fd8c", 
            x"fd18", x"fc08", x"fa04", x"f8f0", 
            x"f9bf", x"fb29", x"fba3", x"fb4c", 
            x"fb9d", x"fdf9", x"02e4", x"09af", 
            x"0faa", x"11ba", x"0fee", x"0dac", 
            x"0d20", x"0d70", x"0d93", x"0dfb", 
            x"0ed6", x"0ecf", x"0bc6", x"05a3", 
            x"001c", x"fea9", x"ffbc", x"ff89", 
            x"fd21", x"fa38", x"f8db", x"f9cf", 
            x"fbf6", x"fe0b", x"0035", x"01fd", 
            x"00b8", x"fafd", x"f4d1", x"f4c0", 
            x"fbf3", x"03ef", x"05de", x"01a1", 
            x"fc9d", x"fb4b", x"fd04", x"fe28", 
            x"fdb5", x"fe54", x"014b", x"0420", 
            x"054e", x"065b", x"07c4", x"07c4", 
            x"06d9", x"086a", x"0cb6", x"0f6d", 
            x"0de6", x"0ad9", x"09a7", x"0953", 
            x"06fb", x"0313", x"0008", x"fde8", 
            x"fb7e", x"f9f4", x"faf6", x"fd58", 
            x"feed", x"febb", x"fc71", x"f8b9", 
            x"f5a7", x"f503", x"f66b", x"f847", 
            x"f978", x"f9d3", x"f98d", x"f8e6", 
            x"f836", x"f84b", x"f9a7", x"fb60", 
            x"fc06", x"fb15", x"f91e", x"f7a4", 
            x"f83b", x"fa8d", x"fc2e", x"fb1e", 
            x"f7d6", x"f4d5", x"f4e4", x"f873", 
            x"fc69", x"fd22", x"fb12", x"fa04", 
            x"fbef", x"fea6", x"ff17", x"fccc", 
            x"f9e9", x"f929", x"fb12", x"fce5", 
            x"fbe3", x"f8dd", x"f6b9", x"f6ba", 
            x"f7d3", x"f8cf", x"fa1e", x"fcbf", 
            x"ff25", x"fe0c", x"f92b", x"f45c", 
            x"f35a", x"f553", x"f643", x"f47a", 
            x"f26e", x"f2a9", x"f528", x"f8c7", 
            x"fc6d", x"fedd", x"ff60", x"fec2", 
            x"fdf1", x"fcd3", x"fbd2", x"fd0e", 
            x"0192", x"068b", x"07e0", x"0511", 
            x"0135", x"fea9", x"fd5b", x"fd8e", 
            x"0043", x"03d9", x"0430", x"fff2", 
            x"f9e5", x"f52a", x"f3bc", x"f642", 
            x"fac8", x"fcfc", x"fa01", x"f469", 
            x"f22a", x"f5e1", x"fc71", x"00e2", 
            x"00c8", x"fd53", x"f9b1", x"f938", 
            x"fd57", x"03ff", x"0976", x"0b96", 
            x"0ae9", x"09d7", x"0a92", x"0ca1", 
            x"0d6b", x"0abc", x"05a5", x"02e4", 
            x"0607", x"0c1a", x"0fb2", x"1066", 
            x"119c", x"13fb", x"1460", x"10ba", 
            x"0ab3", x"05fe", x"0472", x"045b", 
            x"0373", x"02af", x"044b", x"06c8", 
            x"0648", x"02d9", x"00e2", x"034e", 
            x"0820", x"0bef", x"0dce", x"0e10", 
            x"0c99", x"0a97", x"0a55", x"0b42", 
            x"09fb", x"05af", x"014f", x"ff2f", 
            x"ff0f", x"0024", x"0155", x"004a", 
            x"fc0f", x"f728", x"f4b9", x"f587", 
            x"f863", x"fb43", x"fbbe", x"f9d6", 
            x"f92e", x"fca0", x"0218", x"05a3", 
            x"0645", x"057c", x"04df", x"048e", 
            x"030c", x"ff74", x"fc1b", x"fcbb", 
            x"019b", x"06c9", x"0883", x"06f3", 
            x"049c", x"0342", x"0335", x"0432", 
            x"04d3", x"035f", x"ffed", x"fca0", 
            x"faad", x"f970", x"f930", x"fae8", 
            x"fd34", x"fd06", x"f94c", x"f3cd", 
            x"ef46", x"ed20", x"ec4b", x"ead1", 
            x"e895", x"e6a6", x"e54b", x"e4e5", 
            x"e76d", x"ee8a", x"f87c", x"00ea", 
            x"04c6", x"04d2", x"045f", x"0629", 
            x"0a0b", x"0d70", x"0eb7", x"0f0d", 
            x"1013", x"111a", x"10ed", x"10cd", 
            x"1236", x"1336", x"10b3", x"0b5e", 
            x"070a", x"066f", x"094c", x"0c4f", 
            x"0b44", x"0578", x"feda", x"fbb6", 
            x"fc7d", x"fe62", x"ff73", x"fff8", 
            x"ffe7", x"fe21", x"fb99", x"fb39", 
            x"fd60", x"ff84", x"00d4", x"02aa", 
            x"04cb", x"06af", x"0a0d", x"0ea1", 
            x"0f9f", x"0a53", x"0352", x"00c9", 
            x"0279", x"0306", x"003d", x"fddf", 
            x"ff80", x"0304", x"03a7", x"007d", 
            x"fe3e", x"0129", x"06e6", x"097e", 
            x"0626", x"fe36", x"f515", x"ef30", 
            x"ef3a", x"f339", x"f63c", x"f59b", 
            x"f3dd", x"f56b", x"fac1", x"ffdd", 
            x"0219", x"03a7", x"06f2", x"098f", 
            x"07e0", x"02e9", x"ff74", x"0059", 
            x"03f6", x"0613", x"042c", x"007c", 
            x"ff4f", x"0149", x"026b", x"fed7", 
            x"f6da", x"ee7f", x"ea88", x"ec4d", 
            x"f04e", x"f259", x"f247", x"f241", 
            x"f2f6", x"f31b", x"f1f2", x"efee", 
            x"ed96", x"eb6b", x"ea78", x"eb8b", 
            x"ee9e", x"f2c4", x"f617", x"f65c", 
            x"f2f1", x"eeb7", x"ee0a", x"f0db", 
            x"f265", x"f13f", x"f1b5", x"f5a9", 
            x"f916", x"f9bf", x"fbc8", x"01c1", 
            x"06a1", x"050e", x"ffc1", x"fcf3", 
            x"fd7f", x"fe4b", x"fe82", x"ff73", 
            x"0118", x"0271", x"0396", x"055e", 
            x"0726", x"0743", x"05de", x"049e", 
            x"03a3", x"016f", x"fdca", x"f9d1", 
            x"f714", x"f87c", x"ffb2", x"08a8", 
            x"0cd6", x"0aec", x"067c", x"0213", 
            x"fe56", x"fc3c", x"fbfd", x"fbf4", 
            x"fb89", x"fc20", x"fe4a", x"016d", 
            x"05d9", x"0baa", x"1013", x"0fba", 
            x"0bbb", x"0883", x"0857", x"09f5", 
            x"0c9f", x"1138", x"16ae", x"192d", 
            x"1669", x"103c", x"0a8e", x"07c3", 
            x"0696", x"0404", x"000a", x"fd11", 
            x"fb13", x"f8df", x"f7ab", x"f893", 
            x"f9fa", x"fa47", x"f9be", x"f87e", 
            x"f6f8", x"f7c1", x"fd08", x"03e0", 
            x"06cf", x"0606", x"06cd", x"0a87", 
            x"0d2b", x"0d2e", x"0e1a", x"11a2", 
            x"13f4", x"1236", x"0ef8", x"0d22", 
            x"0c0b", x"09de", x"06a0", x"0497", 
            x"06ab", x"0d2d", x"13b6", x"1497", 
            x"0efb", x"074a", x"0249", x"014b", 
            x"014e", x"ff39", x"fc0c", x"fa8a", 
            x"faa4", x"fa2c", x"f906", x"f9eb", 
            x"fd7b", x"ff75", x"fc28", x"f5af", 
            x"f135", x"f174", x"f5b4", x"fb85", 
            x"006a", x"0382", x"04c6", x"0336", 
            x"ff04", x"fc7c", x"ffb2", x"05f2", 
            x"0909", x"07f3", x"0685", x"0749", 
            x"0a0e", x"0d81", x"0ee4", x"0b99", 
            x"04f3", x"0001", x"0000", x"0212", 
            x"0125", x"fcf6", x"fa20", x"fb95", 
            x"ff53", x"011d", x"fe8e", x"f94e", 
            x"f660", x"f944", x"ff85", x"0344", 
            x"0244", x"0015", x"00f2", x"046f", 
            x"06b9", x"05a1", x"021c", x"fe44", 
            x"fc04", x"fbbd", x"fbd0", x"faba", 
            x"f8a4", x"f6af", x"f619", x"f760", 
            x"f961", x"fa36", x"f998", x"f95b", 
            x"fb32", x"fde2", x"fe4d", x"fc88", 
            x"fcf7", x"01b2", x"0695", x"075e", 
            x"04fb", x"0256", x"0040", x"fe81", 
            x"fce4", x"fb3a", x"fa60", x"fc0a", 
            x"0044", x"0485", x"0658", x"068a", 
            x"07a8", x"0982", x"09e2", x"083f", 
            x"0538", x"012b", x"fd61", x"fbb1", 
            x"fb5c", x"faa5", x"fa44", x"fae3", 
            x"f9cf", x"f4dc", x"efce", x"f028", 
            x"f57a", x"fa58", x"fb30", x"f91e", 
            x"f740", x"f641", x"f3eb", x"ef92", 
            x"ecb3", x"eeec", x"f437", x"f720", 
            x"f66c", x"f5fa", x"f81f", x"fb45", 
            x"fda1", x"febd", x"fe7d", x"fe59", 
            x"00d8", x"0516", x"06d9", x"055e", 
            x"04fe", x"08b6", x"0dc2", x"0f9e", 
            x"0db8", x"0a15", x"0691", x"057a", 
            x"0877", x"0cb3", x"0cbe", x"0838", 
            x"0572", x"089b", x"0d35", x"0ccc", 
            x"085d", x"0582", x"04be", x"017d", 
            x"faff", x"f5ce", x"f446", x"f356", 
            x"f04a", x"ed76", x"ed9c", x"ef04", 
            x"ef13", x"eec4", x"f03d", x"f39b", 
            x"f737", x"f9c6", x"fb85", x"fd4d", 
            x"fef0", x"ffeb", x"00e9", x"0228", 
            x"01f3", x"ffb0", x"fe4e", x"00aa", 
            x"046a", x"044f", x"0030", x"fe1d", 
            x"01d4", x"074c", x"0961", x"094b", 
            x"0b51", x"0f5e", x"10c0", x"0cb5", 
            x"056e", x"fecf", x"fa93", x"f7cc", 
            x"f599", x"f540", x"f7ae", x"fad8", 
            x"fc3a", x"fc4c", x"fdd3", x"0173", 
            x"0368", x"ff64", x"f72f", x"f0f5", 
            x"ef5a", x"f0a4", x"f39c", x"f7e0", 
            x"fb96", x"fca2", x"fbf5", x"fd2e", 
            x"0199", x"0588", x"04f3", x"00dd", 
            x"fe30", x"0008", x"049f", x"0872", 
            x"0ae3", x"0d75", x"1023", x"11eb", 
            x"12c4", x"125c", x"0ff9", x"0ce6", 
            x"0c73", x"106f", x"16d3", x"1b2f", 
            x"1a2e", x"13ff", x"0bc5", x"0512", 
            x"019f", x"00bb", x"007d", x"ffd0", 
            x"ff43", x"fff0", x"0267", x"05d9", 
            x"0797", x"0549", x"0053", x"fcb0", 
            x"fb4c", x"f9b8", x"f753", x"f67c", 
            x"f872", x"fbd6", x"ff45", x"0302", 
            x"07c0", x"0bd5", x"0b84", x"05af", 
            x"fe45", x"f9fe", x"f9b7", x"fbaf", 
            x"fea9", x"024f", x"0632", x"0a0f", 
            x"0ea5", x"1400", x"175b", x"15cc", 
            x"1037", x"09f0", x"05da", x"0501", 
            x"04ec", x"019d", x"fb01", x"f51d", 
            x"f23d", x"f126", x"f018", x"ee43", 
            x"ec00", x"eb0d", x"ecb4", x"ef2c", 
            x"ef66", x"ed59", x"ec4d", x"eed2", 
            x"f409", x"f825", x"f76c", x"f2bf", 
            x"eee9", x"ee7c", x"efe5", x"f0ca", 
            x"f185", x"f535", x"fd5f", x"05fb", 
            x"0938", x"066e", x"02e2", x"042d", 
            x"09a8", x"0cc9", x"09de", x"05dd", 
            x"0701", x"0b09", x"0b09", x"06bc", 
            x"03f2", x"0410", x"0223", x"fc10", 
            x"f767", x"f9cc", x"00ff", x"0588", 
            x"0308", x"fbcd", x"f578", x"f38d", 
            x"f57c", x"f838", x"f87d", x"f572", 
            x"f286", x"f380", x"f704", x"f94d", 
            x"f9a7", x"fa24", x"fbf3", x"fec0", 
            x"01e2", x"042e", x"03c7", x"003a", 
            x"fc6a", x"fbd1", x"fdc6", x"fe71", 
            x"fc74", x"fa98", x"fb94", x"fdd2", 
            x"fd7d", x"f98e", x"f590", x"f5a2", 
            x"f848", x"f79a", x"f255", x"ee72", 
            x"f0b2", x"f6b9", x"fb2e", x"fc25", 
            x"fb5b", x"faa5", x"faa7", x"fba3", 
            x"fd19", x"fd7f", x"fc0e", x"fa30", 
            x"f9e2", x"fb13", x"fc22", x"fcc5", 
            x"fe78", x"01e1", x"053a", x"05f5", 
            x"0434", x"02d1", x"0332", x"0394", 
            x"02ca", x"0269", x"03a8", x"05b8", 
            x"07cc", x"096f", x"098e", x"08c5", 
            x"09a5", x"0c56", x"0e08", x"0c52", 
            x"072b", x"0199", x"ffef", x"0301", 
            x"0729", x"09b1", x"0c1c", x"101d", 
            x"1232", x"0d98", x"04de", x"ff09", 
            x"fd6d", x"fb1e", x"f694", x"f463", 
            x"f7b2", x"fe15", x"0375", x"05fa", 
            x"05f8", x"050d", x"0513", x"06cd", 
            x"09be", x"0d32", x"103f", x"115f", 
            x"1002", x"0db1", x"0ca6", x"0dfc", 
            x"1121", x"143d", x"14b4", x"1125", 
            x"0ca2", x"0b4c", x"0b69", x"08b2", 
            x"04ba", x"03f5", x"05b7", x"05d8", 
            x"038a", x"012c", x"000c", x"ffe2", 
            x"006b", x"00ee", x"00b9", x"009f", 
            x"00b8", x"fe09", x"f748", x"f1b8", 
            x"f347", x"f9e5", x"fda8", x"fa81", 
            x"f4c2", x"f363", x"f89a", x"00ff", 
            x"07e3", x"0b62", x"0cd3", x"0e16", 
            x"0ea5", x"0c8f", x"0842", x"04ce", 
            x"039d", x"03d5", x"04ed", x"067d", 
            x"06ca", x"048e", x"0132", x"ffd9", 
            x"017c", x"02c6", x"ffc8", x"fa18", 
            x"f7c0", x"fae1", x"ff8e", x"02a9", 
            x"0545", x"0767", x"058c", x"fea2", 
            x"f738", x"f33d", x"f158", x"efa9", 
            x"efcf", x"f2e6", x"f649", x"f7c4"
        ),
        -- Block 17
        (
            x"f87f", x"f9e5", x"fb99", x"fcfb", 
            x"fca9", x"f8e2", x"f2f9", x"eee6", 
            x"edf5", x"edff", x"eeb6", x"f236", 
            x"f800", x"fc57", x"fd71", x"fd60", 
            x"fe73", x"00e4", x"040f", x"06f4", 
            x"0757", x"03cd", x"fefe", x"fd04", 
            x"fd8b", x"fd44", x"fbe3", x"fc0d", 
            x"feae", x"01f0", x"03dd", x"03f3", 
            x"02ce", x"0135", x"ff26", x"fb92", 
            x"f67c", x"f286", x"f303", x"f8cc", 
            x"00bf", x"05a0", x"03f9", x"fd46", 
            x"f726", x"f651", x"f988", x"fb19", 
            x"f871", x"f5a3", x"f790", x"fd24", 
            x"012e", x"01d1", x"01ed", x"02db", 
            x"0228", x"ff86", x"ff34", x"04b1", 
            x"0d88", x"134a", x"1191", x"0978", 
            x"012c", x"ff5f", x"042b", x"0826", 
            x"054f", x"ff07", x"fd4e", x"025b", 
            x"0925", x"0bfa", x"0920", x"0312", 
            x"feaf", x"fed3", x"0128", x"0095", 
            x"fc62", x"fa9a", x"ff4b", x"0531", 
            x"04cf", x"ffc2", x"fdf2", x"00e7", 
            x"01e4", x"fceb", x"f69b", x"f5d4", 
            x"fc15", x"04ae", x"09b7", x"0951", 
            x"063e", x"034a", x"00a8", x"fe64", 
            x"fdce", x"feff", x"ff95", x"fd80", 
            x"fa6c", x"fa49", x"fdfb", x"0171", 
            x"00e7", x"fd6e", x"f9fa", x"f7b0", 
            x"f6c7", x"f8d7", x"fed1", x"0535", 
            x"0658", x"018f", x"fd43", x"ff39", 
            x"04d6", x"05fd", x"001d", x"f998", 
            x"f81b", x"f98a", x"f993", x"f883", 
            x"f90e", x"fb05", x"fbd3", x"fb0f", 
            x"fb3e", x"fe40", x"030d", x"0757", 
            x"09c2", x"0a19", x"08b6", x"0671", 
            x"03ee", x"01c7", x"0227", x"06f8", 
            x"0d7f", x"1040", x"0ec1", x"0d68", 
            x"0d0d", x"0a30", x"052b", x"039e", 
            x"07a3", x"0b47", x"088f", x"01b7", 
            x"fda9", x"feda", x"01c2", x"026e", 
            x"ffd0", x"fb32", x"f6ea", x"f511", 
            x"f65e", x"f9bb", x"fc11", x"fb11", 
            x"f8cd", x"f90c", x"fb10", x"fae2", 
            x"f82a", x"f6b3", x"f76c", x"f71c", 
            x"f4aa", x"f43a", x"f981", x"010a", 
            x"041c", x"0152", x"fce7", x"fadc", 
            x"fb85", x"fb54", x"f7db", x"f587", 
            x"fac2", x"0612", x"0f0c", x"106e", 
            x"0dd9", x"0de4", x"1199", x"152c", 
            x"15ca", x"136b", x"0fc1", x"0d02", 
            x"0c8e", x"0de1", x"0f59", x"1023", 
            x"10e7", x"126e", x"13ac", x"1365", 
            x"11d3", x"0f28", x"0b1e", x"06d5", 
            x"043a", x"0314", x"009b", x"fbbd", 
            x"f7fd", x"f88c", x"fac1", x"f9ce", 
            x"f62b", x"f3a6", x"f23d", x"ef5b", 
            x"eccd", x"eec2", x"f310", x"f228", 
            x"eabe", x"e5bd", x"ea76", x"f478", 
            x"fa35", x"f970", x"f816", x"fbd8", 
            x"038e", x"0945", x"0a06", x"08da", 
            x"0986", x"0bfc", x"0d71", x"0bcc", 
            x"0948", x"0a8a", x"0fbb", x"1325", 
            x"1093", x"0b72", x"0aa6", x"0e9e", 
            x"103a", x"0b05", x"0293", x"fbc5", 
            x"f67e", x"f1a7", x"eff6", x"f37b", 
            x"f8df", x"fb46", x"fa49", x"f92e", 
            x"fa20", x"fced", x"0084", x"0338", 
            x"02f3", x"fef9", x"f9a0", x"f70f", 
            x"f99c", x"fe7e", x"ff06", x"f90c", 
            x"f35f", x"f52f", x"fc61", x"0152", 
            x"0174", x"00cc", x"02bb", x"05ab", 
            x"066b", x"0403", x"0022", x"fd7c", 
            x"fccd", x"fbb6", x"f765", x"f0e6", 
            x"ecfc", x"edf1", x"f0b3", x"f223", 
            x"f2a5", x"f356", x"f412", x"f4c7", 
            x"f5e1", x"f68b", x"f48d", x"f0a3", 
            x"efa9", x"f447", x"fb5a", x"00c3", 
            x"03f1", x"0735", x"0c26", x"114c", 
            x"139b", x"1109", x"0b30", x"0753", 
            x"09d0", x"10c1", x"14e9", x"11d0", 
            x"0af9", x"06d3", x"06fe", x"08cc", 
            x"0942", x"05bf", x"fe1b", x"f6ae", 
            x"f4c0", x"f805", x"f9ed", x"f52b", 
            x"ebea", x"e501", x"e49c", x"e8f9", 
            x"ecf8", x"ed08", x"ea46", x"e864", 
            x"e92d", x"ead9", x"eb11", x"ea4d", 
            x"eaa4", x"ed6f", x"f290", x"f7c3", 
            x"f99a", x"f8cc", x"fb25", x"028e", 
            x"08b1", x"08ac", x"0682", x"0773", 
            x"0972", x"077a", x"01bf", x"fdb3", 
            x"fe66", x"00dc", x"00cf", x"fdd6", 
            x"fa76", x"f890", x"f79f", x"f69a", 
            x"f621", x"f703", x"f847", x"f841", 
            x"f5ec", x"f157", x"ec75", x"ea24", 
            x"eb49", x"ee64", x"f1fb", x"f59f", 
            x"f924", x"fd6b", x"03f1", x"0ae2", 
            x"0c8b", x"0691", x"fe5c", x"fa81", 
            x"fb74", x"fe81", x"0348", x"0a0c", 
            x"0fab", x"106e", x"0dd4", x"0bf1", 
            x"0b07", x"0964", x"0801", x"08db", 
            x"0bd4", x"0ed9", x"0ed2", x"0a5c", 
            x"041f", x"00c0", x"0211", x"04ab", 
            x"03a1", x"fe88", x"fa7a", x"fc05", 
            x"012c", x"04bb", x"0565", x"0570", 
            x"054d", x"0284", x"fc84", x"f783", 
            x"f7fb", x"fc6c", x"ffc5", x"002b", 
            x"ff40", x"ff34", x"0228", x"0866", 
            x"0e96", x"10f0", x"0fbf", x"0e45", 
            x"0d7a", x"0b84", x"0862", x"06d1", 
            x"079b", x"08b6", x"091a", x"093d", 
            x"0807", x"054c", x"05d3", x"0c86", 
            x"12f0", x"1117", x"0941", x"044b", 
            x"0498", x"0473", x"fff6", x"fa12", 
            x"f791", x"f925", x"fbc1", x"fce2", 
            x"fc44", x"fa8f", x"f841", x"f5bd", 
            x"f3da", x"f3e7", x"f661", x"fa9e", 
            x"ffc5", x"04e4", x"0839", x"092b", 
            x"0a35", x"0cf2", x"0dd9", x"08cc", 
            x"006c", x"fbe7", x"fde0", x"018f", 
            x"01d1", x"ffa8", x"fffe", x"04d7", 
            x"0a70", x"0b61", x"071b", x"0270", 
            x"00f2", x"01bd", x"0320", x"0411", 
            x"02df", x"ffc1", x"fe76", x"00ff", 
            x"03d3", x"038c", x"0258", x"02e3", 
            x"038f", x"020f", x"fdb0", x"f6ee", 
            x"f0fb", x"eff8", x"f2e6", x"f3f4", 
            x"f152", x"f032", x"f4f7", x"fc84", 
            x"0048", x"fdf1", x"f831", x"f281", 
            x"ef45", x"f01a", x"f4cb", x"fa81", 
            x"fe90", x"0181", x"0490", x"05a8", 
            x"0288", x"fddd", x"fbff", x"fc78", 
            x"fb76", x"f8e9", x"f8d2", x"fb9f", 
            x"fcd6", x"fb39", x"fb0c", x"ff43", 
            x"05bc", x"0aca", x"0c3c", x"097c", 
            x"03b8", x"feb3", x"fe22", x"fff3", 
            x"fe80", x"f9a5", x"f699", x"f6a7", 
            x"f690", x"f5bc", x"f68d", x"f885", 
            x"f7ec", x"f3e4", x"f1bd", x"f726", 
            x"01a0", x"08df", x"09ac", x"082c", 
            x"07be", x"072f", x"04ed", x"0256", 
            x"0187", x"01f9", x"01c8", x"00f3", 
            x"017b", x"0514", x"0a88", x"0da5", 
            x"0b24", x"048d", x"fe63", x"fa70", 
            x"f779", x"f570", x"f5e9", x"f9c1", 
            x"00ca", x"08ce", x"0cd0", x"0a10", 
            x"0449", x"0198", x"031c", x"0446", 
            x"01fd", x"fe8e", x"fdd9", x"00f6", 
            x"05a1", x"0953", x"0c60", x"1036", 
            x"1421", x"16cc", x"187b", x"1964", 
            x"1775", x"10ba", x"0873", x"04b3", 
            x"0672", x"08d4", x"0a0d", x"0d69", 
            x"1355", x"16bb", x"1475", x"0f7e", 
            x"0c46", x"0be7", x"0bad", x"0895", 
            x"0389", x"0196", x"05ce", x"0bdf", 
            x"0cb5", x"0834", x"0618", x"0aed", 
            x"10b6", x"0f60", x"0790", x"0054", 
            x"fdf7", x"fe2a", x"fcdb", x"fa14", 
            x"f850", x"f81a", x"f85b", x"f9a7", 
            x"fe7f", x"0743", x"1071", x"15a5", 
            x"1594", x"12c6", x"114f", x"124a", 
            x"11af", x"0b64", x"020e", x"fd0d", 
            x"ff08", x"0425", x"0873", x"0a65", 
            x"08c6", x"044b", x"0123", x"01a4", 
            x"0231", x"feb1", x"f9eb", x"f962", 
            x"fba1", x"fa13", x"f3de", x"ef8d", 
            x"f0cd", x"f3e8", x"f520", x"f5f3", 
            x"f8ae", x"fc87", x"004c", x"0407", 
            x"069e", x"04c5", x"fc73", x"f175", 
            x"ecb3", x"f28a", x"fb97", x"fd8e", 
            x"f8cd", x"f5dc", x"f890", x"fd2d", 
            x"ff0c", x"fc75", x"f752", x"f3d2", 
            x"f4a7", x"f8a3", x"fd23", x"0107", 
            x"0368", x"02c4", x"ff92", x"fc43", 
            x"f9b2", x"f6d3", x"f39b", x"f119", 
            x"f000", x"f165", x"f656", x"fcd3", 
            x"ffe7", x"fed7", x"fe72", x"0074", 
            x"0136", x"ff0d", x"fc73", x"fb98", 
            x"fc56", x"fe15", x"0074", x"01b6", 
            x"0073", x"ff32", x"0227", x"08e7", 
            x"0e88", x"0f04", x"09f1", x"02df", 
            x"ff67", x"0170", x"0432", x"01b6", 
            x"faa0", x"f501", x"f45e", x"f6b6", 
            x"f8af", x"f86d", x"f60d", x"f3df", 
            x"f46a", x"f6ae", x"f69a", x"f319", 
            x"efcf", x"eef6", x"ef2b", x"eff2", 
            x"f241", x"f527", x"f70a", x"f984", 
            x"fef5", x"04eb", x"0614", x"02dd", 
            x"01da", x"05be", x"09e3", x"09ba", 
            x"05ee", x"02b1", x"0310", x"0521", 
            x"0526", x"0323", x"01b7", x"017b", 
            x"00bf", x"fe83", x"fbe2", x"fa6f", 
            x"fa94", x"fc51", x"fed8", x"ffe5", 
            x"feaa", x"fd11", x"fc53", x"fc70", 
            x"fdc7", x"fee4", x"fc1b", x"f4f7", 
            x"ee48", x"ec8b", x"ef0b", x"f1f4", 
            x"f315", x"f342", x"f4d1", x"f9f9", 
            x"01af", x"062c", x"0324", x"fced", 
            x"fa86", x"fb8d", x"fb02", x"f952", 
            x"fb81", x"002a", x"0040", x"fc3a", 
            x"fc31", x"00da", x"0236", x"fc7a", 
            x"f4f9", x"f2b4", x"f6cf", x"fcc3", 
            x"005c", x"0203", x"034c", x"033f", 
            x"0130", x"ff7c", x"ffb8", x"0072", 
            x"009f", x"012d", x"020b", x"0156", 
            x"ff68", x"0097", x"07af", x"1089", 
            x"13e1", x"1002", x"09ca", x"06bb", 
            x"07d0", x"08c7", x"0645", x"0357", 
            x"0424", x"060c", x"041b", x"0030", 
            x"0016", x"04b9", x"09b2", x"0b19", 
            x"0859", x"034b", x"ff42", x"ff21", 
            x"011b", x"ffe7", x"fb32", x"f841", 
            x"f8dd", x"f9fb", x"faf7", x"fdfc", 
            x"01ff", x"0357", x"0112", x"fd47", 
            x"fb22", x"fd56", x"02a4", x"0548", 
            x"0222", x"fe24", x"ff0e", x"0217", 
            x"0048", x"f934", x"f374", x"f423", 
            x"fa06", x"ffad", x"ffd0", x"fa9d", 
            x"f777", x"fd4a", x"082c", x"0c14", 
            x"0417", x"f8b5", x"f3ae", x"f535", 
            x"f8a8", x"fca7", x"01e6", x"06cc", 
            x"092f", x"0a14", x"0aee", x"0a02", 
            x"064b", x"042b", x"07d2", x"0d12", 
            x"0b80", x"0243", x"fa14", x"fa8a", 
            x"0134", x"071c", x"0a25", x"0ac3", 
            x"0753", x"002f", x"fabe", x"faf3", 
            x"fe2e", x"0003", x"006b", x"014f", 
            x"0189", x"ff24", x"fbaa", x"fb10", 
            x"fed5", x"0355", x"02b9", x"fb34", 
            x"f223", x"efda", x"f6b4", x"0054", 
            x"05ee", x"06e1", x"0547", x"0254", 
            x"002b", x"013c", x"0527", x"0910", 
            x"0b1c", x"0bcd", x"0ae4", x"06b9", 
            x"00f8", x"feef", x"017c", x"0301", 
            x"002f", x"fbe9", x"fa14", x"fbdd", 
            x"ff60", x"00bc", x"fe19", x"fa92", 
            x"fb29", x"005b", x"04ab", x"0339", 
            x"fe18", x"fc0c", x"0005", x"0584", 
            x"06a4", x"0289", x"fc88", x"f8fd", 
            x"fa49", x"fdec", x"ff8a", x"fee6", 
            x"fe75", x"feda", x"ff63", x"ffed", 
            x"008a", x"00f7", x"0044", x"fcc7", 
            x"f6fe", x"f3c2", x"f6dd", x"fcef", 
            x"ffbe", x"fe18", x"fbb4", x"fb3e", 
            x"fb1e", x"f818", x"f201", x"ed0d", 
            x"ede3", x"f3e7", x"fa69", x"fecf", 
            x"0137", x"00d1", x"fce5", x"f8f4", 
            x"fa2f", x"ffde", x"02fb", x"005a", 
            x"fdce", x"0161", x"087d", x"0c61", 
            x"0b72", x"093d", x"08d0", x"0a13", 
            x"0af2", x"0a21", x"085d", x"071b", 
            x"074b", x"098f", x"0d2a", x"0f2a", 
            x"0d2d", x"08c3", x"0607", x"0776", 
            x"0c0e", x"1025", x"102e", x"0c46", 
            x"0968", x"0c12", x"1101", x"10a3", 
            x"09b2", x"0215", x"fe1f", x"fd2b", 
            x"fdae", x"fe36", x"fc57", x"f824"
        ),
        -- Block 16
        (
            x"f5db", x"f7d7", x"fb04", x"fba9", 
            x"f9b6", x"f742", x"f5bf", x"f522", 
            x"f5b5", x"f8e6", x"fee4", x"0577", 
            x"0967", x"093a", x"07ab", x"0880", 
            x"0bbf", x"0f22", x"10c7", x"0f8e", 
            x"0bfa", x"0847", x"057b", x"032f", 
            x"02f0", x"05f7", x"0874", x"0597", 
            x"ffdd", x"fe02", x"00dc", x"0314", 
            x"00bc", x"fa42", x"f31d", x"efcc", 
            x"f1b1", x"f4ed", x"f4bb", x"f166", 
            x"efb2", x"f277", x"f6f7", x"f911", 
            x"f7eb", x"f542", x"f318", x"f275", 
            x"f2fa", x"f42c", x"f77e", x"fe34", 
            x"062a", x"0b71", x"0b82", x"06e7", 
            x"01e1", x"006a", x"00bc", x"ff20", 
            x"fd32", x"ff1b", x"0373", x"04c1", 
            x"0224", x"fff9", x"ff67", x"fd3e", 
            x"f8a8", x"f496", x"f231", x"ef83", 
            x"eceb", x"edc9", x"f211", x"f508", 
            x"f33b", x"ed7c", x"e7d5", x"e74d", 
            x"edc5", x"f7a8", x"fe90", x"ff78", 
            x"fdb6", x"fdac", x"ff9a", x"0248", 
            x"05de", x"0a1b", x"0d7e", x"0efa", 
            x"0f7d", x"106e", x"104b", x"0bf3", 
            x"0394", x"fbf6", x"fa22", x"fd0f", 
            x"fe90", x"fc73", x"faae", x"fba5", 
            x"fc97", x"fb75", x"f9ce", x"f949", 
            x"fa9a", x"fecd", x"04fd", x"082e", 
            x"0419", x"fba6", x"f650", x"f73f", 
            x"fa1f", x"fb31", x"fdd0", x"0551", 
            x"0d19", x"0f91", x"0eab", x"0f19", 
            x"109c", x"1062", x"0e90", x"0da4", 
            x"0dd5", x"0d0f", x"0b49", x"0ab9", 
            x"0b87", x"0ad7", x"077d", x"03fc", 
            x"0175", x"fe2d", x"fba0", x"fd69", 
            x"0114", x"01a9", x"0055", x"0155", 
            x"03cf", x"0364", x"ff03", x"f98d", 
            x"f606", x"f666", x"fc04", x"04e1", 
            x"0b89", x"0ca9", x"0b99", x"0db7", 
            x"1247", x"14d5", x"14d0", x"1495", 
            x"151b", x"161d", x"1682", x"13c1", 
            x"0d09", x"06d9", x"062f", x"08ec", 
            x"0856", x"01e9", x"fa03", x"f65a", 
            x"f80f", x"fc21", x"fed1", x"fda8", 
            x"fa73", x"fa0b", x"fcd6", x"fd7b", 
            x"f926", x"f4c3", x"f6bb", x"fdbf", 
            x"0341", x"046f", x"0319", x"0155", 
            x"00b6", x"01ba", x"0288", x"0175", 
            x"ff09", x"fc11", x"f975", x"fa18", 
            x"0000", x"0862", x"0e27", x"0ef5", 
            x"0c34", x"0957", x"0928", x"0b5e", 
            x"0cf2", x"0b35", x"06f8", x"0481", 
            x"05e4", x"0758", x"0539", x"01a1", 
            x"000c", x"008d", x"0183", x"016a", 
            x"fed5", x"fa5c", x"f7cb", x"fa67", 
            x"006c", x"0436", x"0228", x"fcbe", 
            x"f93e", x"f959", x"fb31", x"fd25", 
            x"fda6", x"facb", x"f5b0", x"f293", 
            x"f2f7", x"f379", x"f1e8", x"f1b1", 
            x"f5e1", x"fab4", x"fa9e", x"f76a", 
            x"f72f", x"faa3", x"fdac", x"fecd", 
            x"ff4f", x"fe06", x"f962", x"f403", 
            x"f2b6", x"f79b", x"ffca", x"049b", 
            x"0112", x"f7db", x"f162", x"f1ef", 
            x"f5fb", x"f89d", x"f87a", x"f59c", 
            x"f0e1", x"ee17", x"f064", x"f4a5", 
            x"f52a", x"f208", x"f036", x"f1d5", 
            x"f481", x"f693", x"f7a3", x"f625", 
            x"f315", x"f33b", x"f7ed", x"fc5f", 
            x"fc23", x"f8b0", x"f6cf", x"f7f6", 
            x"fa06", x"fbdf", x"fde0", x"0006", 
            x"019a", x"01e7", x"0196", x"025b", 
            x"049d", x"0667", x"0699", x"06bd", 
            x"06e6", x"049e", x"00ed", x"0055", 
            x"0304", x"0417", x"00d3", x"fb48", 
            x"f66d", x"f3f3", x"f55f", x"fb4d", 
            x"01f9", x"0375", x"ff14", x"faa3", 
            x"fac0", x"fd95", x"fe0e", x"f9be", 
            x"f366", x"f06b", x"f344", x"f8e0", 
            x"fc9b", x"fd2c", x"fc6c", x"fb7d", 
            x"f934", x"f63a", x"f6d7", x"fbd3", 
            x"fedf", x"fb0b", x"f3e0", x"f17f", 
            x"f775", x"00c4", x"0629", x"0652", 
            x"044f", x"01b9", x"fff5", x"023a", 
            x"084b", x"0ba2", x"0656", x"fb53", 
            x"f3fb", x"f48b", x"f7ea", x"f989", 
            x"fb6d", x"fe5b", x"fdd6", x"f896", 
            x"f547", x"f96f", x"0005", x"ffe8", 
            x"f938", x"f421", x"f4e6", x"f914", 
            x"fde0", x"02bd", x"0711", x"09f1", 
            x"0b4e", x"0b7a", x"09aa", x"0535", 
            x"ff82", x"fc0a", x"fe1b", x"04da", 
            x"0b1b", x"0d9d", x"0e1c", x"0ea8", 
            x"0e3a", x"0b21", x"05f8", x"0148", 
            x"ffd4", x"02ac", x"0879", x"0e70", 
            x"11c5", x"1001", x"0989", x"046f", 
            x"06a4", x"0d97", x"1158", x"0e40", 
            x"0702", x"0011", x"fc18", x"fbcb", 
            x"fe5a", x"0096", x"ff90", x"fd40", 
            x"fdf8", x"0143", x"0297", x"0060", 
            x"fe0d", x"fd4c", x"fb58", x"f820", 
            x"f79c", x"faab", x"fe6a", x"0182", 
            x"03df", x"03a6", x"00b2", x"febc", 
            x"ff83", x"fff7", x"fdf7", x"fc37", 
            x"fe2d", x"03b1", x"0a60", x"1014", 
            x"12c4", x"116d", x"0d97", x"095a", 
            x"0515", x"0053", x"fb79", x"f8dc", 
            x"fbb0", x"03c3", x"0ba7", x"0d87", 
            x"095d", x"04f0", x"043e", x"044a", 
            x"00f1", x"fb57", x"f832", x"fb52", 
            x"0331", x"08b1", x"07b7", x"0502", 
            x"05e5", x"08a7", x"094d", x"080a", 
            x"0795", x"06fb", x"02cf", x"fd68", 
            x"fd64", x"0259", x"04ba", x"02b0", 
            x"02ea", x"0873", x"0cd4", x"0b13", 
            x"0831", x"097c", x"0bae", x"0abc", 
            x"0870", x"06db", x"0547", x"0444", 
            x"05d2", x"097e", x"0ccf", x"0de2", 
            x"0bdd", x"0791", x"045c", x"0542", 
            x"0824", x"074a", x"0192", x"fc3e", 
            x"faa2", x"f9f1", x"f793", x"f53d", 
            x"f50e", x"f791", x"fca3", x"0223", 
            x"03fc", x"00c2", x"fb95", x"f74e", 
            x"f3b0", x"f0ca", x"f027", x"f191", 
            x"f3f8", x"f7de", x"fd39", x"0241", 
            x"0605", x"0807", x"06bd", x"0211", 
            x"fc9e", x"f853", x"f57f", x"f5e9", 
            x"fb20", x"01e2", x"0580", x"060c", 
            x"05cd", x"0455", x"0185", x"0152", 
            x"05be", x"08a6", x"0356", x"f8ff", 
            x"f16e", x"ee62", x"edb9", x"efa2", 
            x"f3b2", x"f648", x"f514", x"f17f", 
            x"ed6f", x"e9ad", x"e766", x"e8d1", 
            x"ee27", x"f350", x"f558", x"f71a", 
            x"fc4f", x"0360", x"06e8", x"0596", 
            x"0414", x"050a", x"05ca", x"04f6", 
            x"04f1", x"067f", x"08a6", x"0c69", 
            x"119b", x"1378", x"0fb5", x"0b91", 
            x"0aec", x"09c4", x"0549", x"030a", 
            x"07a6", x"0d1b", x"0ade", x"03a1", 
            x"00cd", x"03d1", x"0634", x"040e", 
            x"ff13", x"fa79", x"f81c", x"f755", 
            x"f58a", x"f24b", x"f20f", x"f7ac", 
            x"fd09", x"fa89", x"f40e", x"f413", 
            x"fb61", x"0047", x"fde5", x"fa74", 
            x"fd17", x"04ab", x"0ac4", x"0b1e", 
            x"0777", x"065b", x"0bd2", x"130b", 
            x"1304", x"0a3d", x"01ad", x"0245", 
            x"0a69", x"1098", x"0e3b", x"0542", 
            x"fcf3", x"fad9", x"fdc3", x"ffb3", 
            x"fd50", x"f968", x"f7d1", x"f7ae", 
            x"f6ab", x"f690", x"fa0a", x"0041", 
            x"078c", x"0f13", x"142b", x"133c", 
            x"0d2e", x"0867", x"092c", x"0c64", 
            x"0c7b", x"092b", x"0764", x"094c", 
            x"0b49", x"0a6d", x"07ed", x"04b5", 
            x"00ac", x"fec9", x"01bf", x"0627", 
            x"05e4", x"0060", x"fb20", x"faa3", 
            x"fced", x"fcd8", x"f9a8", x"f713", 
            x"f6b5", x"f6f4", x"f777", x"f93c", 
            x"fbc3", x"fd3a", x"fd15", x"fd00", 
            x"fdf2", x"fee3", x"ff17", x"ff8f", 
            x"0100", x"021a", x"0106", x"fe48", 
            x"fc1e", x"fb46", x"fb46", x"fc3a", 
            x"fc4b", x"f8d8", x"f4ad", x"f59c", 
            x"faf6", x"fdd3", x"fc50", x"fca5", 
            x"00ac", x"0057", x"f7e8", x"effe", 
            x"ef6f", x"f12d", x"ef8e", x"ed3c", 
            x"ed65", x"edb6", x"ed35", x"f01c", 
            x"f854", x"002e", x"0112", x"fc75", 
            x"fa60", x"fe7c", x"030d", x"02be", 
            x"00fe", x"0365", x"08a8", x"0a77", 
            x"06be", x"030a", x"0445", x"06fe", 
            x"061e", x"0437", x"068e", x"0b8f", 
            x"0d76", x"0b00", x"07c0", x"0555", 
            x"01c0", x"fcbe", x"f9b1", x"f9c9", 
            x"f925", x"f6a8", x"f7a5", x"fe9a", 
            x"059c", x"0660", x"012e", x"fa90", 
            x"f684", x"f5e4", x"f778", x"faba", 
            x"fe9a", x"ff6f", x"fba3", x"f818", 
            x"faf0", x"01d9", x"035e", x"fcab", 
            x"f72e", x"fb61", x"03c2", x"04d0", 
            x"fd8c", x"f806", x"fa73", x"ff52", 
            x"0010", x"fe8a", x"fe7c", x"fff2", 
            x"02a0", x"064a", x"07ff", x"0542", 
            x"00cf", x"ff7d", x"00d9", x"0114", 
            x"fffc", x"ffe3", x"012f", x"02f6", 
            x"052d", x"0873", x"0ae2", x"087d", 
            x"02e8", x"004e", x"0080", x"fe8a", 
            x"fa95", x"f875", x"f863", x"f838", 
            x"f7fd", x"f944", x"fc6e", x"0019", 
            x"011e", x"fc68", x"f43c", x"f0bb", 
            x"f5d8", x"fc0a", x"fae8", x"f69b", 
            x"f83d", x"fd87", x"fd11", x"f6a5", 
            x"f1bb", x"f0a0", x"f0f1", x"f2c0", 
            x"f6ad", x"f9d4", x"fa7c", x"fbbe", 
            x"ffa7", x"0346", x"0481", x"05b4", 
            x"0889", x"0a1c", x"07f0", x"0603", 
            x"08dc", x"0c68", x"0a70", x"04e5", 
            x"0182", x"0119", x"0098", x"febd", 
            x"fdfa", x"ffd2", x"0136", x"fe52", 
            x"f77a", x"f1c8", x"f22c", x"f73d", 
            x"fb05", x"fb04", x"f975", x"f89a", 
            x"f84a", x"f775", x"f6c1", x"f885", 
            x"fdeb", x"054a", x"0b56", x"0ddd", 
            x"0d93", x"0c9d", x"0b5b", x"084f", 
            x"042c", x"026b", x"0427", x"05df", 
            x"05ef", x"08c7", x"103a", x"1633", 
            x"15cb", x"1109", x"0b96", x"06f5", 
            x"03ab", x"01e3", x"00ff", x"00d0", 
            x"0159", x"0057", x"faf7", x"f3fe", 
            x"f3c7", x"fd47", x"06be", x"056a", 
            x"fce2", x"f9bf", x"fff1", x"072a", 
            x"07a4", x"02be", x"fe88", x"fec7", 
            x"02e8", x"07a2", x"0acf", x"0c33", 
            x"0b65", x"0876", x"0585", x"0583", 
            x"0a33", x"115e", x"145f", x"0e7b", 
            x"03fe", x"ff79", x"0525", x"0bc5", 
            x"07ee", x"fc67", x"f6fa", x"fda2", 
            x"0751", x"091d", x"0264", x"fa5d", 
            x"f7a0", x"f9a7", x"f995", x"f394", 
            x"ed87", x"f022", x"fa5c", x"025c", 
            x"01ef", x"fd1d", x"fbbc", x"ff1a", 
            x"0078", x"fbda", x"f73b", x"f9fb", 
            x"02f2", x"0ac5", x"0d4d", x"0e8f", 
            x"13cb", x"1a34", x"1c18", x"1a7b", 
            x"19ba", x"19bf", x"1821", x"1578", 
            x"13b4", x"12d2", x"1263", x"12bf", 
            x"126e", x"0e38", x"05f8", x"fd78", 
            x"f8ae", x"f99a", x"fe98", x"01f8", 
            x"fefb", x"f7c8", x"f3fb", x"f6da", 
            x"fb0d", x"fb6d", x"fa24", x"fb6d", 
            x"003e", x"06a7", x"0ba2", x"0ce3", 
            x"0a36", x"06d0", x"0725", x"0a25", 
            x"0a35", x"065a", x"024f", x"0050", 
            x"006f", x"0253", x"0603", x"0b8c", 
            x"0f56", x"0b5b", x"0058", x"f66e", 
            x"f202", x"ef89", x"ec43", x"eba7", 
            x"f0b6", x"f7c1", x"fb64", x"fd5c", 
            x"030b", x"0a78", x"0bbe", x"0481", 
            x"f9a0", x"f007", x"eaf4", x"ec99", 
            x"f25e", x"f625", x"f690", x"f7ee", 
            x"fc2d", x"ff51", x"fe11", x"fb99", 
            x"fbe2", x"fcc3", x"fab2", x"f736", 
            x"f567", x"f4c6", x"f42d", x"f514", 
            x"f7da", x"fa6b", x"fbe3", x"fd68", 
            x"ff9e", x"018d", x"0294", x"02d2", 
            x"01a1", x"ff69", x"ff7a", x"034b", 
            x"0681", x"046e", x"ffa7", x"fda3", 
            x"fe88", x"ff82", x"0018", x"00be", 
            x"0072", x"fd93", x"f718", x"ef53", 
            x"ec8e", x"f0c6", x"f45a", x"f050", 
            x"e8fd", x"e712", x"ea7c", x"ebce", 
            x"e799", x"e1e6", x"e01d", x"e2d6", 
            x"e56a", x"e40f", x"e24b", x"e5e6", 
            x"ebaa", x"eb48", x"e681", x"e689"
        ),
        -- Block 15
        (
            x"eb4f", x"ecbd", x"e9f3", x"ea20", 
            x"efda", x"f55d", x"f76d", x"f981", 
            x"fc71", x"fc44", x"f97e", x"fa6f", 
            x"00f1", x"0697", x"05bb", x"010f", 
            x"ff81", x"02ae", x"054f", x"042c", 
            x"02be", x"03f1", x"04c1", x"01f4", 
            x"fe07", x"fd18", x"fe5c", x"fefa", 
            x"feec", x"fe5c", x"fcb8", x"fc41", 
            x"fe30", x"fe58", x"fb80", x"fb83", 
            x"0010", x"0163", x"fad2", x"f2c1", 
            x"f13d", x"f598", x"f992", x"fa35", 
            x"f925", x"f8d1", x"fac3", x"fd58", 
            x"fc5a", x"f8df", x"f9de", x"00a3", 
            x"074f", x"0add", x"0c2c", x"0b55", 
            x"0a05", x"0bec", x"0fe6", x"0f77", 
            x"08b6", x"024a", x"0290", x"07f4", 
            x"0c99", x"0e5b", x"0f91", x"11b1", 
            x"1348", x"128f", x"0ee9", x"0874", 
            x"017b", x"fdfb", x"fdd3", x"fcb3", 
            x"fa80", x"fc7a", x"04e9", x"0fca", 
            x"1697", x"1558", x"0f6a", x"0cf9", 
            x"10bf", x"1582", x"161f", x"1310", 
            x"10b9", x"1180", x"1207", x"0d2b", 
            x"03cd", x"fda0", x"ffc3", x"069a", 
            x"0bc3", x"0cc0", x"09db", x"0600", 
            x"0722", x"0ddd", x"113f", x"0bf7", 
            x"05a8", x"066d", x"0a1d", x"0799", 
            x"fd3f", x"f25c", x"f092", x"fa20", 
            x"0679", x"0b39", x"0697", x"012c", 
            x"055a", x"115d", x"1807", x"12b1", 
            x"08a4", x"0383", x"055b", x"09bb", 
            x"0b8c", x"0976", x"0559", x"0102", 
            x"fce6", x"fa16", x"fa94", x"fdf9", 
            x"0068", x"00b7", x"02b6", x"07b6", 
            x"0abd", x"06d7", x"fe0a", x"f81d", 
            x"fa3c", x"ffeb", x"ff55", x"f6b0", 
            x"efa3", x"f152", x"f668", x"f5e2", 
            x"efac", x"eb5f", x"ece2", x"f060", 
            x"f212", x"f245", x"f136", x"ef37", 
            x"f0ad", x"f8f1", x"02b7", x"0749", 
            x"0877", x"0901", x"05e8", x"ff8b", 
            x"fc91", x"ff02", x"00b8", x"fdc6", 
            x"fb53", x"ffaf", x"0853", x"0d80", 
            x"0b89", x"05b4", x"01af", x"0106", 
            x"009d", x"fe3e", x"fb97", x"fc44", 
            x"01c2", x"0946", x"0f31", x"10d0", 
            x"0b53", x"0090", x"f93f", x"fb20", 
            x"025c", x"083c", x"0baf", x"0fd8", 
            x"1440", x"1498", x"1121", x"0f25", 
            x"0f63", x"0cbe", x"058a", x"fed3", 
            x"fc1d", x"fbb5", x"fcc7", x"0030", 
            x"046f", x"069b", x"0652", x"0514", 
            x"040f", x"045f", x"06c6", x"09a6", 
            x"0b05", x"0d25", x"11b1", x"13d3", 
            x"0f5b", x"0842", x"05ad", x"0818", 
            x"0838", x"02a9", x"fe07", x"ff78", 
            x"04fb", x"0c89", x"1334", x"127f", 
            x"0a2a", x"0331", x"0290", x"0333", 
            x"00d1", x"fed3", x"ffa3", x"ff6c", 
            x"fcbe", x"fbad", x"fc68", x"fa2b", 
            x"f55a", x"f3a8", x"f5e0", x"f78f", 
            x"f920", x"fe0d", x"0188", x"fcb7", 
            x"f5ae", x"f5c8", x"f8a9", x"f532", 
            x"edd2", x"eadb", x"ecb3", x"ee9b", 
            x"f014", x"f22f", x"f241", x"ef17", 
            x"ee57", x"f5e9", x"023c", x"08c3", 
            x"050a", x"fe49", x"fce7", x"ffa6", 
            x"ffec", x"fbe8", x"f6d7", x"f3de", 
            x"f48a", x"f8ef", x"fe74", x"019a", 
            x"025b", x"031b", x"03a5", x"0217", 
            x"00d1", x"04df", x"0cda", x"112b", 
            x"0f6f", x"0d12", x"0b90", x"0676", 
            x"fe1f", x"f7c7", x"f608", x"f7c2", 
            x"f8f2", x"f4b7", x"ec60", x"e91c", 
            x"f0ca", x"fbf6", x"fe18", x"f611", 
            x"eccf", x"e6c3", x"e362", x"e63f", 
            x"f1b4", x"fca1", x"fc0b", x"f37e", 
            x"ef9a", x"f3be", x"f7e6", x"f61d", 
            x"f15f", x"f04e", x"f4f3", x"fa89", 
            x"fc89", x"fccd", x"ff37", x"03ad", 
            x"07bd", x"0b3b", x"0f49", x"1167", 
            x"0d21", x"0495", x"00bd", x"0511", 
            x"0b43", x"0ea0", x"11d2", x"16e2", 
            x"1a35", x"1763", x"0fbe", x"0a3f", 
            x"09c2", x"0744", x"fd0c", x"f155", 
            x"ed96", x"f2aa", x"faea", x"0000", 
            x"fdf9", x"f6aa", x"ef80", x"ea71", 
            x"e6f1", x"e6cf", x"ea7a", x"ee0d", 
            x"ee12", x"ec14", x"edbb", x"f5bf", 
            x"fdbc", x"fd92", x"f774", x"f3f4", 
            x"f579", x"f7b3", x"f742", x"f5f6", 
            x"f85c", x"fe5d", x"0262", x"03aa", 
            x"0764", x"0c6b", x"0b22", x"03f8", 
            x"00e3", x"058b", x"0ad3", x"0b8b", 
            x"0a4c", x"09bd", x"087f", x"0719", 
            x"0868", x"09aa", x"055e", x"fd9e", 
            x"f862", x"f613", x"f4d7", x"f634", 
            x"faa3", x"fe30", x"fe61", x"fe6b", 
            x"0145", x"04b1", x"067e", x"07d5", 
            x"08f6", x"0873", x"06bb", x"04f6", 
            x"015f", x"fb24", x"f726", x"fabb", 
            x"0305", x"0816", x"0742", x"0521", 
            x"05a5", x"066e", x"044b", x"0163", 
            x"006f", x"0080", x"00c4", x"0157", 
            x"0193", x"01ab", x"016a", x"fe87", 
            x"f9a3", x"f81b", x"fa97", x"f93d", 
            x"f030", x"e94c", x"f04b", x"007e", 
            x"0903", x"020f", x"f44d", x"ec6a", 
            x"f041", x"fc19", x"0545", x"0448", 
            x"fcf2", x"f861", x"fbe1", x"069b", 
            x"11c5", x"1515", x"0f96", x"091a", 
            x"08c9", x"0ca2", x"0dea", x"0bfe", 
            x"0b9e", x"0c54", x"0979", x"04ea", 
            x"0459", x"0812", x"0c8a", x"0fad", 
            x"1154", x"1225", x"1180", x"0de2", 
            x"08a9", x"05e7", x"06b8", x"0714", 
            x"0384", x"febe", x"fda5", x"ffbe", 
            x"005b", x"fe1e", x"fb1e", x"f75a", 
            x"f2e5", x"f176", x"f4f1", x"f998", 
            x"fb2f", x"f8ad", x"f3ce", x"f0ea", 
            x"f2e2", x"f5a6", x"f38f", x"ef74", 
            x"f0f1", x"f7f3", x"fd21", x"fe7f", 
            x"0154", x"06f6", x"0a55", x"0a99", 
            x"0d4b", x"1346", x"15a5", x"10ee", 
            x"0aa0", x"0919", x"0c41", x"0f05", 
            x"0ebc", x"0fb5", x"15c8", x"1b98", 
            x"19a2", x"1150", x"0b2f", x"0c37", 
            x"0fa3", x"0d42", x"0512", x"0018", 
            x"052c", x"114f", x"1bef", x"1fa7", 
            x"1d0d", x"186a", x"1524", x"11bd", 
            x"0b77", x"0535", x"0434", x"0691", 
            x"0467", x"fbec", x"f5bb", x"f8d9", 
            x"001c", x"0156", x"fb23", x"f4a1", 
            x"f270", x"f2bf", x"f0a1", x"e90a", 
            x"df3b", x"db30", x"dfdb", x"e617", 
            x"e6d2", x"e575", x"e957", x"f165", 
            x"f6e3", x"f8e2", x"fbb5", x"feb7", 
            x"fd80", x"f9cf", x"f9db", x"fe4f", 
            x"01c9", x"019a", x"01b7", x"066a", 
            x"0ce7", x"0df8", x"084a", x"0389", 
            x"0619", x"0c48", x"0c38", x"016b", 
            x"f46a", x"f131", x"f7f7", x"fe9a", 
            x"fd78", x"f59c", x"ef43", x"f21d", 
            x"fb6e", x"00c0", x"fda9", x"f853", 
            x"f736", x"f8a9", x"f869", x"f766", 
            x"f8c3", x"fc0d", x"fea4", x"ff0b", 
            x"fdf3", x"fd9d", x"ff7f", x"0200", 
            x"01c4", x"0001", x"03b9", x"0e8a", 
            x"16d6", x"1468", x"0a74", x"0029", 
            x"f870", x"f37a", x"f1a4", x"f2ec", 
            x"f660", x"f9d4", x"faaa", x"f835", 
            x"f51f", x"f526", x"f8a3", x"fac5", 
            x"f798", x"f2b4", x"f309", x"f99e", 
            x"00af", x"01e3", x"fd9b", x"fbca", 
            x"0131", x"0874", x"0acf", x"0959", 
            x"09ab", x"0d12", x"0ebe", x"0b40", 
            x"059e", x"03a8", x"08d4", x"1210", 
            x"160d", x"101d", x"0790", x"0634", 
            x"0c76", x"1226", x"10dd", x"0b45", 
            x"07e1", x"082f", x"089d", x"06bc", 
            x"041d", x"01ee", x"fd91", x"f5fb", 
            x"f0d4", x"f4f0", x"003b", x"08aa", 
            x"081e", x"0276", x"fdfc", x"fb9c", 
            x"f8ea", x"f5ac", x"f4b3", x"f82b", 
            x"fdee", x"00cc", x"ff4f", x"fd5b", 
            x"fea8", x"03cc", x"0a4d", x"0cee", 
            x"079c", x"fd37", x"f61f", x"f715", 
            x"fc3f", x"ffe2", x"021b", x"0515", 
            x"066e", x"039f", x"0009", x"ff7c", 
            x"001f", x"feff", x"fd34", x"fd3a", 
            x"fee6", x"001e", x"008f", x"0329", 
            x"094f", x"0ec6", x"0d1e", x"0332", 
            x"faa2", x"ffbf", x"0fe4", x"198e", 
            x"1216", x"02ac", x"fbac", x"ff70", 
            x"0264", x"ffbc", x"ff54", x"0306", 
            x"01b6", x"f92f", x"f2bb", x"f344", 
            x"f523", x"f251", x"eb76", x"e5ce", 
            x"e5c8", x"ead4", x"ef20", x"ed63", 
            x"e7a6", x"e52d", x"e845", x"ebea", 
            x"eccb", x"ed89", x"f05b", x"f2e5", 
            x"f26d", x"ef35", x"ec90", x"ef0c", 
            x"f679", x"fde8", x"039d", x"0a58", 
            x"12be", x"177d", x"12fd", x"082f", 
            x"ffca", x"fcdb", x"faf8", x"f7a9", 
            x"f613", x"f82d", x"fb45", x"fd09", 
            x"fdab", x"fc4a", x"f803", x"f449", 
            x"f54e", x"fa1c", x"ff62", x"043d", 
            x"08d4", x"0c48", x"0d09", x"0a7b", 
            x"07cd", x"089d", x"0abd", x"098d", 
            x"051f", x"01b3", x"02d2", x"07d7", 
            x"0d21", x"10b3", x"1233", x"1026", 
            x"0a48", x"0516", x"049a", x"0496", 
            x"ff54", x"f878", x"f70e", x"fa98", 
            x"fdc1", x"fdc1", x"f9d0", x"f21b", 
            x"eba5", x"ecdb", x"f3fc", x"f993", 
            x"fbc5", x"0027", x"087d", x"0ca3", 
            x"072b", x"ffd0", x"ff43", x"0286", 
            x"02b8", x"00ae", x"0142", x"03c6", 
            x"044d", x"0408", x"067f", x"0965", 
            x"081a", x"04b6", x"0545", x"09c4", 
            x"0cae", x"0ba7", x"0871", x"0442", 
            x"00b9", x"0121", x"0456", x"03ff", 
            x"fed6", x"facf", x"faba", x"fabe", 
            x"f8d5", x"f8aa", x"fc9d", x"01d3", 
            x"05c2", x"085a", x"0814", x"037e", 
            x"fe70", x"fd3d", x"fd82", x"fb65", 
            x"f898", x"f782", x"f63c", x"f464", 
            x"f648", x"fda6", x"0586", x"09b0", 
            x"0bf6", x"0e37", x"0dc3", x"07e6", 
            x"fe61", x"f596", x"f017", x"edcc", 
            x"ef5f", x"f5a3", x"fdbb", x"0442", 
            x"0b0d", x"13a3", x"185a", x"13c5", 
            x"0afd", x"0823", x"0c22", x"0eb2", 
            x"0d10", x"0db0", x"12f3", x"15f9", 
            x"12a9", x"0e36", x"0db9", x"0f23", 
            x"0db2", x"0830", x"00b4", x"fa4b", 
            x"f899", x"fd33", x"038e", x"0491", 
            x"fe2c", x"f435", x"eca1", x"eaf3", 
            x"ecf5", x"ee81", x"ef80", x"f21f", 
            x"f600", x"f8aa", x"f958", x"fab0", 
            x"ff62", x"047c", x"03d6", x"fe06", 
            x"fb63", x"0080", x"079b", x"098b", 
            x"0712", x"0522", x"07c8", x"0f8b", 
            x"149f", x"0ddf", x"ff9b", x"f794", 
            x"fb6f", x"03ce", x"0793", x"0633", 
            x"049e", x"04fe", x"06d4", x"09a8", 
            x"0b71", x"0a56", x"093b", x"0c3d", 
            x"1117", x"11de", x"0d2f", x"06c8", 
            x"0280", x"020a", x"03f0", x"0295", 
            x"faca", x"f282", x"f17a", x"f6f8", 
            x"fc5c", x"fe1b", x"fdd7", x"fe0f", 
            x"0016", x"03e8", x"07cd", x"0819", 
            x"00d5", x"f292", x"e528", x"e105", 
            x"e55d", x"e9cb", x"e996", x"e97f", 
            x"ef5a", x"f805", x"fce0", x"fde5", 
            x"ff40", x"0280", x"0603", x"067a", 
            x"019e", x"fa48", x"f7ff", x"fe53", 
            x"0687", x"0931", x"082a", x"07c4", 
            x"0663", x"0140", x"fbe0", x"fc5b", 
            x"0152", x"02ea", x"fe1d", x"f8c6", 
            x"f953", x"fd83", x"fc35", x"f1e4", 
            x"e5ab", x"df25", x"ddf8", x"de78", 
            x"e047", x"e4ba", x"eaf0", x"ef18", 
            x"edc4", x"e7d4", x"e27e", x"e3db", 
            x"ebbe", x"f18a", x"ef6b", x"ea90", 
            x"ea95", x"eef4", x"f202", x"f394", 
            x"fa4e", x"0681", x"0cd5", x"067f", 
            x"fbd5", x"f7b6", x"fa99", x"fefc", 
            x"01db", x"0209", x"fcbf", x"f1cf", 
            x"e877", x"e834", x"ee9c", x"f2ff", 
            x"f202", x"ef03", x"ed26", x"ec8b", 
            x"ec5e", x"edbb", x"f2dd", x"f970", 
            x"fb58", x"f7d8", x"f4bc", x"f597", 
            x"f963", x"feaa", x"031e", x"03be", 
            x"00c7", x"fef7", x"0197", x"065d", 
            x"0a4d", x"0e1d", x"1265", x"1451"
        ),
        -- Block 14
        (
            x"12d5", x"1182", x"128f", x"1351", 
            x"11b7", x"0fc8", x"0fb0", x"0fb8", 
            x"0d82", x"0a9b", x"0a1c", x"0ce4", 
            x"10df", x"12a4", x"1192", x"10f0", 
            x"121e", x"10e1", x"0a85", x"049e", 
            x"05ed", x"0c4e", x"1090", x"103d", 
            x"0dc9", x"0a84", x"0629", x"00fe", 
            x"fbc2", x"f85e", x"f85b", x"fa12", 
            x"facd", x"fb0c", x"fd42", x"013c", 
            x"04f8", x"0904", x"0db7", x"10fc", 
            x"12d7", x"153b", x"170f", x"15b4", 
            x"13b9", x"1764", x"1f00", x"2013", 
            x"1856", x"1265", x"14d3", x"19fe", 
            x"1ab2", x"16c2", x"124c", x"10ed", 
            x"132b", x"1452", x"0f7b", x"08c7", 
            x"088d", x"0dcb", x"0fa6", x"0bdc", 
            x"083e", x"0602", x"010a", x"facc", 
            x"f9a9", x"fe10", x"0136", x"fdc3", 
            x"f5ff", x"f22b", x"f74b", x"00d5", 
            x"071b", x"0765", x"03e9", x"00e2", 
            x"01a8", x"073e", x"0e44", x"0e9e", 
            x"0537", x"fc1d", x"fe7e", x"07d3", 
            x"0adc", x"04e8", x"fd53", x"f801", 
            x"f550", x"f877", x"0196", x"0794", 
            x"02ac", x"fa17", x"fb77", x"06d6", 
            x"0f41", x"0d0e", x"04a9", x"fec7", 
            x"ff25", x"0127", x"ff8d", x"fd3c", 
            x"fee4", x"01cd", x"011a", x"fdb3", 
            x"fb26", x"fa83", x"fbdf", x"ff76", 
            x"0303", x"03da", x"02ee", x"023f", 
            x"00a6", x"fb6f", x"f276", x"e8e1", 
            x"e2db", x"e39a", x"e985", x"ecc9", 
            x"e8f2", x"e6e9", x"f04e", x"fcf8", 
            x"fdb4", x"f3a2", x"ed3e", x"f1ce", 
            x"fb2c", x"fefc", x"fa04", x"f477", 
            x"f840", x"054c", x"122f", x"14aa", 
            x"0acb", x"fe89", x"fba9", x"0264", 
            x"0ac8", x"1061", x"1318", x"12da", 
            x"1014", x"0b76", x"0536", x"ff7e", 
            x"fb66", x"f5ca", x"eeeb", x"ef72", 
            x"fc03", x"08cb", x"06c0", x"f7ef", 
            x"ea87", x"e5ae", x"e4af", x"e239", 
            x"e006", x"e237", x"e9a2", x"f3f6", 
            x"fb73", x"fad6", x"f68f", x"f865", 
            x"008b", x"05ca", x"0275", x"fa36", 
            x"f474", x"f58a", x"fd64", x"0844", 
            x"0f8f", x"0f51", x"0bb7", x"0b4a", 
            x"0e80", x"11cf", x"134c", x"1243", 
            x"0e47", x"0849", x"01c0", x"fbea", 
            x"f88a", x"f945", x"fd45", x"ffb6", 
            x"fbb9", x"f41a", x"f148", x"f585", 
            x"fb17", x"fe00", x"0017", x"0306", 
            x"0317", x"fdd4", x"f84c", x"f5bf", 
            x"f182", x"ebdb", x"ee67", x"fa36", 
            x"02b2", x"009a", x"fc38", x"0093", 
            x"0c0f", x"1218", x"0b47", x"ff4b", 
            x"fb4c", x"0257", x"0c9b", x"1228", 
            x"111b", x"0d91", x"0d7a", x"1005", 
            x"0da8", x"041f", x"fa60", x"f7b1", 
            x"fc40", x"020f", x"0450", x"0387", 
            x"0291", x"0359", x"0601", x"07e0", 
            x"0469", x"fbbc", x"f584", x"f6f8", 
            x"fabd", x"f970", x"f3eb", x"eff2", 
            x"f12f", x"f835", x"021a", x"0883", 
            x"07f2", x"04fb", x"06b5", x"0d52", 
            x"1105", x"0c8a", x"0494", x"0093", 
            x"019d", x"03d8", x"03e8", x"0114", 
            x"fd2f", x"fb90", x"ff52", x"075b", 
            x"0d3f", x"0c6a", x"07cd", x"04a3", 
            x"02e2", x"fec9", x"f80c", x"f1ef", 
            x"ecd4", x"e71a", x"e316", x"e53f", 
            x"ee00", x"f758", x"fa4f", x"f7a4", 
            x"f6b6", x"fab6", x"fec7", x"fec3", 
            x"fb09", x"f4db", x"f035", x"f25a", 
            x"f9d8", x"0018", x"02db", x"0365", 
            x"00e6", x"fc3e", x"fb60", x"0316", 
            x"0f43", x"14df", x"0d7e", x"ff50", 
            x"f690", x"f86f", x"fdd4", x"fb96", 
            x"f0b7", x"e913", x"eea3", x"fbcd", 
            x"02f9", x"00a7", x"fc0b", x"f95e", 
            x"f7ba", x"f891", x"fbd3", x"faf6", 
            x"f38b", x"ee43", x"f24a", x"fa01", 
            x"fb9f", x"f7ff", x"f899", x"00bc", 
            x"094d", x"0b8e", x"099c", x"08df", 
            x"08a6", x"044a", x"fcda", x"fb3b", 
            x"02d9", x"098c", x"0615", x"fde3", 
            x"fb37", x"fe17", x"00cf", x"02b7", 
            x"050f", x"0363", x"fa83", x"f2a3", 
            x"f4de", x"fb9b", x"fcbe", x"fab8", 
            x"fcf4", x"021e", x"0448", x"020a", 
            x"fe4c", x"fd6f", x"02ad", x"0bcd", 
            x"119b", x"10ee", x"0e64", x"0e8d", 
            x"1093", x"1161", x"0ea0", x"0879", 
            x"0305", x"02a1", x"05a0", x"04c2", 
            x"fefc", x"fecf", x"0a81", x"17a2", 
            x"1827", x"0ced", x"02a5", x"01e5", 
            x"079f", x"0a32", x"049f", x"fd63", 
            x"fe78", x"0790", x"0f14", x"0fcf", 
            x"0d8f", x"0bea", x"097e", x"0771", 
            x"0b26", x"1324", x"15ab", x"0edd", 
            x"068d", x"0542", x"0a39", x"0e7d", 
            x"0f20", x"0eaa", x"0d7e", x"09ff", 
            x"0682", x"05a1", x"050d", x"0082", 
            x"f7d3", x"f13d", x"f334", x"fb91", 
            x"01eb", x"03d5", x"0764", x"0f6d", 
            x"1607", x"160b", x"10fb", x"099b", 
            x"01f2", x"fcc0", x"fc05", x"fed8", 
            x"0165", x"025d", x"060c", x"0d07", 
            x"109b", x"0ea6", x"0d68", x"1051", 
            x"1133", x"099b", x"fe99", x"fa05", 
            x"fbc2", x"fc89", x"f9e5", x"f585", 
            x"ef56", x"e751", x"e0bc", x"e053", 
            x"e5d3", x"eb22", x"ede4", x"f044", 
            x"f07a", x"ed50", x"ed1b", x"f454", 
            x"fce0", x"fee1", x"fa64", x"f430", 
            x"efd8", x"ef15", x"f222", x"f7f4", 
            x"fea4", x"0403", x"06ff", x"06ad", 
            x"0216", x"fdbf", x"00fd", x"0934", 
            x"0b44", x"03ea", x"fada", x"f6f6", 
            x"f7e3", x"f907", x"f758", x"f3f2", 
            x"f1cd", x"f0ef", x"edff", x"e84c", 
            x"e485", x"e7a0", x"efdf", x"f61a", 
            x"f80b", x"fab6", x"ff52", x"ff34", 
            x"f66e", x"eb1b", x"e711", x"ece2", 
            x"f566", x"f993", x"fb4a", x"ffb4", 
            x"0534", x"0620", x"03aa", x"04ac", 
            x"095a", x"09d3", x"02d2", x"faf8", 
            x"f7ea", x"f836", x"fc78", x"067c", 
            x"0ec8", x"0d45", x"066a", x"034b", 
            x"0672", x"0c62", x"0e3d", x"068f", 
            x"f91b", x"f194", x"f57f", x"fb36", 
            x"f63f", x"ead7", x"e905", x"f32e", 
            x"fb97", x"fbc4", x"fab6", x"fdf9", 
            x"0357", x"05da", x"01e2", x"f81c", 
            x"ee5f", x"e9dd", x"eb27", x"f05f", 
            x"f66c", x"fa8f", x"fe75", x"0499", 
            x"09b8", x"0921", x"042a", x"0113", 
            x"0425", x"0b14", x"0fff", x"0feb", 
            x"0d76", x"0daf", x"1285", x"1844", 
            x"1964", x"14a7", x"106a", x"1453", 
            x"1d5d", x"1f12", x"1399", x"0291", 
            x"f6ff", x"f5a4", x"fb02", x"fd8b", 
            x"f7dd", x"f042", x"ef8c", x"f677", 
            x"ffa5", x"04f2", x"034e", x"fe34", 
            x"fb1d", x"fa1a", x"f94e", x"fa9a", 
            x"fe82", x"ff6d", x"f8ac", x"f0ff", 
            x"f4fd", x"042f", x"10d4", x"146f", 
            x"13d5", x"10c0", x"0997", x"031d", 
            x"0400", x"0a53", x"0dbf", x"0a28", 
            x"033e", x"fdb7", x"f948", x"f4f8", 
            x"f569", x"ff5b", x"0c92", x"0ee7", 
            x"01d5", x"f07f", x"e74b", x"e7bc", 
            x"ebe0", x"ef77", x"f0db", x"eec6", 
            x"eb4a", x"ead9", x"ef5c", x"f71f", 
            x"feb0", x"01a5", x"fc06", x"f004", 
            x"e7dc", x"eb8f", x"f79a", x"01c3", 
            x"0464", x"012d", x"fcbe", x"fb48", 
            x"fdec", x"02b7", x"06cf", x"0880", 
            x"09cc", x"0da8", x"1147", x"0ed3", 
            x"06e7", x"00aa", x"0053", x"01ec", 
            x"ff4c", x"f9e8", x"f894", x"fae6", 
            x"f88e", x"f0eb", x"ee8c", x"f529", 
            x"faad", x"f929", x"f6b4", x"f83a", 
            x"fc0d", x"fdf2", x"fa3a", x"f4f8", 
            x"f822", x"022a", x"05b4", x"feed", 
            x"f7fd", x"f877", x"fdee", x"02c5", 
            x"0486", x"04bc", x"0524", x"0560", 
            x"04b3", x"0364", x"035a", x"084d", 
            x"12b0", x"1ae3", x"19ee", x"13fb", 
            x"1249", x"15b5", x"16da", x"1022", 
            x"029b", x"f6cf", x"f6a5", x"fee8", 
            x"0180", x"fa24", x"f3c8", x"f81e", 
            x"02e4", x"0927", x"06df", x"01ad", 
            x"0093", x"0270", x"ffff", x"f733", 
            x"ef81", x"efba", x"f4f0", x"f837", 
            x"f9c5", x"ff03", x"08cf", x"12d4", 
            x"1986", x"1b5a", x"199a", x"1817", 
            x"16fc", x"11f9", x"08e6", x"00d0", 
            x"fd51", x"fe87", x"0220", x"05ed", 
            x"0a80", x"0f37", x"0f5e", x"0987", 
            x"0325", x"ffb2", x"faf9", x"f16f", 
            x"e94f", x"eb6e", x"f4df", x"f90e", 
            x"f337", x"ecfb", x"eeff", x"f493", 
            x"f505", x"f0df", x"ef2c", x"f295", 
            x"f7f0", x"fc4d", x"fe9a", x"fde7", 
            x"fba7", x"fc24", x"0112", x"067f", 
            x"0683", x"001e", x"fa34", x"fc8a", 
            x"0518", x"0a0b", x"0605", x"fe6d", 
            x"fd19", x"0504", x"0e3d", x"0f99", 
            x"0925", x"02f5", x"03a4", x"08eb", 
            x"0ba9", x"0a46", x"09f8", x"0d21", 
            x"0e41", x"088e", x"000c", x"fba7", 
            x"fc81", x"0088", x"05e1", x"094a", 
            x"08c3", x"0786", x"0948", x"0ad0", 
            x"050c", x"f882", x"eeb2", x"ed12", 
            x"ef8c", x"f16a", x"f26c", x"f3d8", 
            x"f600", x"f9cb", x"00d5", x"08d7", 
            x"0c11", x"09ce", x"079f", x"07e9", 
            x"0876", x"08c5", x"0942", x"08c2", 
            x"0852", x"09d7", x"0c38", x"0fd2", 
            x"16d5", x"1edc", x"22e9", x"221f", 
            x"1e1f", x"18cb", x"15ad", x"155e", 
            x"145d", x"1256", x"11e9", x"12c5", 
            x"1397", x"15c6", x"19a8", x"198f", 
            x"0f8f", x"ffdd", x"f629", x"f6a2", 
            x"f796", x"f04a", x"e75c", x"e756", 
            x"ed92", x"f10b", x"f109", x"f153", 
            x"efd2", x"e992", x"e44c", x"e615", 
            x"ea3a", x"ec96", x"f41c", x"035c", 
            x"0d74", x"086f", x"fc1b", x"f62f", 
            x"f954", x"fddc", x"ff10", x"fef5", 
            x"ffa1", x"01d3", x"056b", x"0759", 
            x"069c", x"06fb", x"0927", x"0814", 
            x"ffeb", x"f5d7", x"f5df", x"023a", 
            x"0d12", x"0b81", x"0404", x"01bd", 
            x"049a", x"06d9", x"08fa", x"0d44", 
            x"0f3a", x"0a44", x"02ee", x"fff7", 
            x"00d0", x"00bb", x"fc36", x"f377", 
            x"ebda", x"ebe8", x"f401", x"fdaa", 
            x"03aa", x"06ae", x"080c", x"05cc", 
            x"fe2c", x"f456", x"edb2", x"eb25", 
            x"ea88", x"ec9c", x"f1ef", x"f655", 
            x"f603", x"f1ce", x"ec94", x"ea28", 
            x"edc7", x"f425", x"f439", x"eb6a", 
            x"e525", x"ebca", x"f6bc", x"f77a", 
            x"f029", x"ed14", x"f2aa", x"fc30", 
            x"01ed", x"0000", x"fb2c", x"fa52", 
            x"fda7", x"0113", x"0122", x"fda3", 
            x"fabd", x"fd01", x"0515", x"0f4d", 
            x"171c", x"1b37", x"1c5d", x"1b65", 
            x"1abe", x"1b72", x"19b3", x"12fa", 
            x"0afc", x"06e2", x"0848", x"0c49", 
            x"0da4", x"0a58", x"0401", x"fe0a", 
            x"ff3b", x"0a47", x"14ae", x"11d7", 
            x"0418", x"f83c", x"f483", x"f39d", 
            x"ef13", x"e8fc", x"e64b", x"e5be", 
            x"e4f6", x"e5b3", x"e9c0", x"efdf", 
            x"f658", x"fc05", x"fe6c", x"fb76", 
            x"f56c", x"f24e", x"f5b1", x"fc10", 
            x"ffd8", x"00eb", x"032c", x"0803", 
            x"0ca5", x"0d76", x"0999", x"0505", 
            x"0562", x"099b", x"0ba9", x"09a6", 
            x"063f", x"0280", x"fc45", x"f3fc", 
            x"ef3e", x"f007", x"f1d3", x"f34f", 
            x"f7e8", x"febe", x"02cc", x"02d2", 
            x"01bb", x"0211", x"01fd", x"fd69", 
            x"f563", x"f0d1", x"f445", x"f9f3", 
            x"f6c4", x"ebab", x"e6a1", x"ed6c", 
            x"f43f", x"f055", x"e8b1", x"eb09", 
            x"f696", x"fe15", x"fb53", x"f3f8", 
            x"edb4", x"e9e8", x"eb43", x"f34b", 
            x"fbcd", x"fe27", x"fe16", x"0341", 
            x"0c22", x"10dd", x"0fb8", x"0cf1", 
            x"0954", x"040e", x"ffce", x"fed3", 
            x"0168", x"07ab", x"0e72", x"1141", 
            x"1081", x"0f39", x"0f6c", x"11b0"
        ),
        -- Block 13
        (
            x"11fc", x"0afe", x"00ab", x"fd39", 
            x"01b7", x"0562", x"03da", x"003b", 
            x"fe7d", x"0042", x"052b", x"0b81", 
            x"0eee", x"0b79", x"0412", x"ff96", 
            x"ffbb", x"022e", x"0559", x"0792", 
            x"0758", x"063f", x"067c", x"065e", 
            x"0372", x"ff61", x"fd7b", x"fdb9", 
            x"ff99", x"04d4", x"0c11", x"103b", 
            x"1007", x"0ed0", x"0db0", x"0ac3", 
            x"072b", x"05f0", x"0728", x"08f3", 
            x"08d5", x"05d5", x"0445", x"0a31", 
            x"16da", x"21c7", x"21c0", x"17e8", 
            x"1183", x"1561", x"1934", x"143f", 
            x"0be0", x"0720", x"06e8", x"09ce", 
            x"0d67", x"0dbb", x"0727", x"fcac", 
            x"f754", x"fa5d", x"ffa9", x"0143", 
            x"fe04", x"f780", x"f2bd", x"f693", 
            x"0182", x"06d8", x"0067", x"f933", 
            x"fae7", x"ffe6", x"ff85", x"fae8", 
            x"fa31", x"009f", x"081a", x"0b29", 
            x"09cf", x"0343", x"f91c", x"f3e2", 
            x"f80c", x"fded", x"fe47", x"ff18", 
            x"080c", x"117a", x"0f9b", x"06d4", 
            x"03ae", x"07d6", x"0a6e", x"066e", 
            x"0181", x"00a0", x"00a2", x"001c", 
            x"0180", x"03fe", x"055b", x"043e", 
            x"fde9", x"f2c5", x"eba0", x"ef0a", 
            x"f521", x"f3cd", x"edfc", x"ec76", 
            x"f2f1", x"fe19", x"0596", x"0416", 
            x"fec0", x"fdc1", x"ffec", x"fe10", 
            x"f730", x"f218", x"f2ee", x"f3d6", 
            x"f061", x"ef4a", x"f4ab", x"f905", 
            x"f6b4", x"f041", x"e8a8", x"e32f", 
            x"e57a", x"efd5", x"f7a9", x"f1c9", 
            x"e20e", x"d920", x"de43", x"e5bf", 
            x"e4bf", x"e0a1", x"e26d", x"e9c8", 
            x"efec", x"eef3", x"ea44", x"ecfb", 
            x"f7af", x"fb12", x"efd6", x"e430", 
            x"e4ef", x"eb33", x"ed21", x"eece", 
            x"f6ce", x"006e", x"02ba", x"fcbd", 
            x"f5e0", x"f2f8", x"f187", x"f1d2", 
            x"f7c6", x"ff8e", x"0136", x"fe30", 
            x"fe4a", x"049a", x"0e18", x"14da", 
            x"1546", x"11df", x"0d12", x"0564", 
            x"fd73", x"fc5a", x"0220", x"091d", 
            x"0db7", x"0d5b", x"08b5", x"06ca", 
            x"0b73", x"1051", x"0ee4", x"08d4", 
            x"0147", x"f70c", x"ecca", x"ec76", 
            x"f744", x"ff36", x"fb8f", x"f49d", 
            x"f375", x"f4bb", x"f1ec", x"ed7c", 
            x"ef92", x"f9c8", x"0367", x"039e", 
            x"fb7d", x"f491", x"f729", x"00cb", 
            x"0642", x"0181", x"f947", x"f904", 
            x"038c", x"10f6", x"17cb", x"145f", 
            x"0a01", x"0143", x"0218", x"0c45", 
            x"161a", x"1510", x"0b07", x"066f", 
            x"0e4d", x"1690", x"133a", x"0a41", 
            x"05b8", x"03e3", x"0141", x"023e", 
            x"096c", x"105d", x"1126", x"1031", 
            x"14f1", x"1cd9", x"1f96", x"1ae5", 
            x"127a", x"0b4f", x"095d", x"0bfd", 
            x"0d7b", x"0b9d", x"0d14", x"1737", 
            x"21b6", x"209b", x"1602", x"0d51", 
            x"0b0c", x"08d3", x"00ba", x"f7d2", 
            x"f696", x"f9ed", x"f7b4", x"ef7c", 
            x"ea70", x"ed7a", x"f38f", x"f57a", 
            x"f395", x"f2f9", x"f4ef", x"f753", 
            x"f836", x"f822", x"fad0", x"00eb", 
            x"0416", x"00f8", x"fde5", x"0005", 
            x"0309", x"03b5", x"07a2", x"1080", 
            x"181f", x"1bd9", x"1b46", x"147d", 
            x"0b9c", x"0918", x"0c62", x"0c1e", 
            x"0623", x"02f3", x"05d5", x"0769", 
            x"035e", x"ff5f", x"0145", x"057a", 
            x"047c", x"fe70", x"fa6f", x"fc27", 
            x"014c", x"05b8", x"04f3", x"ff5b", 
            x"fc93", x"0039", x"0377", x"02d7", 
            x"0381", x"05a0", x"06de", x"0c51", 
            x"16c1", x"1abe", x"11e4", x"0507", 
            x"ffb6", x"0456", x"0bf5", x"0f65", 
            x"0f61", x"0e74", x"0c76", x"0ce7", 
            x"1400", x"1b4d", x"16df", x"083a", 
            x"fe0f", x"fd5d", x"fc98", x"f842", 
            x"f719", x"fab3", x"fc59", x"f803", 
            x"f379", x"f74a", x"0145", x"06be", 
            x"02d8", x"fa1a", x"f3f6", x"f50f", 
            x"fc2e", x"0263", x"020f", x"fdc9", 
            x"fca9", x"0114", x"0633", x"057e", 
            x"fda7", x"f536", x"f602", x"0252", 
            x"1048", x"15a6", x"13c3", x"123f", 
            x"11e0", x"0b86", x"fd4e", x"ef6b", 
            x"e967", x"e9bf", x"ea1a", x"e818", 
            x"e629", x"e67d", x"e87a", x"eae6", 
            x"edc6", x"ef6e", x"edab", x"eb31", 
            x"eb7d", x"ebbb", x"e954", x"e84f", 
            x"e987", x"e67d", x"dcb0", x"d3f2", 
            x"d459", x"db0f", x"df6a", x"e008", 
            x"e253", x"e793", x"eaa5", x"e92c", 
            x"e8da", x"ef7f", x"fbfe", x"0633", 
            x"0468", x"f9ea", x"f730", x"00e3", 
            x"083f", x"0455", x"fce4", x"fa7f", 
            x"fd50", x"0000", x"fd86", x"f798", 
            x"f2e2", x"ef16", x"eaff", x"e97c", 
            x"ebff", x"efbe", x"f2e0", x"f533", 
            x"f4c0", x"f124", x"f0e9", x"f888", 
            x"ff8d", x"fcfd", x"f5a6", x"f13a", 
            x"f129", x"f5e6", x"fc9a", x"ffa2", 
            x"00c1", x"060d", x"0f13", x"15e3", 
            x"17d7", x"1986", x"1ece", x"2189", 
            x"1b8d", x"12ec", x"10bf", x"142d", 
            x"14e2", x"0d82", x"017c", x"f9a5", 
            x"fc4f", x"0616", x"0a67", x"040b", 
            x"fef2", x"03bc", x"06ac", x"fdc4", 
            x"f390", x"f569", x"ffed", x"0678", 
            x"03bb", x"fd02", x"fc3f", x"06d3", 
            x"1526", x"1672", x"05b8", x"f43c", 
            x"f407", x"0390", x"1382", x"16b3", 
            x"0f16", x"0abd", x"10c2", x"1a25", 
            x"1e50", x"1b43", x"146e", x"0fab", 
            x"10c7", x"1537", x"15db", x"1073", 
            x"0c7a", x"116b", x"1ad0", x"1d70", 
            x"172c", x"1212", x"13a2", x"1113", 
            x"02fc", x"f65c", x"f677", x"fa94", 
            x"f83b", x"f56b", x"fbcb", x"05fb", 
            x"07ac", x"fee8", x"f2d1", x"ea57", 
            x"e8d4", x"ece0", x"f211", x"f5f1", 
            x"fa1c", x"ffc9", x"023d", x"fd51", 
            x"f6f2", x"f7b6", x"fed7", x"0454", 
            x"0428", x"0385", x"0780", x"0c6c", 
            x"0cec", x"08f2", x"04b0", x"058e", 
            x"0d6c", x"179b", x"1dc4", x"1e5f", 
            x"1aa5", x"1360", x"0b50", x"0773", 
            x"08ae", x"0995", x"0540", x"fe81", 
            x"fd99", x"0362", x"03ee", x"f88d", 
            x"ecc9", x"eb6b", x"ed7d", x"e8d4", 
            x"e24f", x"e5ee", x"f1a7", x"f55c", 
            x"ecc8", x"e6b0", x"edde", x"fb93", 
            x"0279", x"fde5", x"f5ae", x"f4b6", 
            x"fc7b", x"0500", x"06c2", x"02d2", 
            x"fe8e", x"fcec", x"00a9", x"0cbc", 
            x"1dae", x"2774", x"217a", x"1406", 
            x"0e6d", x"0fef", x"0bda", x"00fd", 
            x"f7f6", x"f320", x"f077", x"f1b7", 
            x"f847", x"fc86", x"f4af", x"e5bc", 
            x"deb6", x"e231", x"e615", x"e7f0", 
            x"ec83", x"f19c", x"f1e8", x"ee7b", 
            x"eccf", x"ef33", x"f153", x"ef38", 
            x"ecde", x"f067", x"f94d", x"0209", 
            x"0557", x"0551", x"091e", x"0e19", 
            x"0b73", x"03d8", x"0041", x"012a", 
            x"0229", x"00e9", x"fe37", x"fca2", 
            x"fb4f", x"f7e7", x"f54e", x"f7f4", 
            x"fe0f", x"00d0", x"fcfe", x"f7e8", 
            x"f993", x"0080", x"01c9", x"fae2", 
            x"f69e", x"f9f8", x"fd26", x"fc16", 
            x"fd35", x"0409", x"09af", x"0895", 
            x"03ce", x"fd67", x"f65e", x"f779", 
            x"04ea", x"11d5", x"123e", x"0b49", 
            x"083f", x"0c5e", x"128e", x"13c6", 
            x"0dec", x"068f", x"0405", x"067a", 
            x"08ab", x"0627", x"0152", x"ff70", 
            x"ffc5", x"fd27", x"f5d4", x"ee93", 
            x"ef4e", x"f849", x"fd11", x"f540", 
            x"ebd1", x"eef1", x"f9b0", x"feb0", 
            x"fd52", x"ff00", x"0741", x"1002", 
            x"13c2", x"1284", x"0ea0", x"0bec", 
            x"0ddd", x"1146", x"10cc", x"1019", 
            x"135e", x"12d1", x"06f2", x"f6e8", 
            x"f062", x"f4d1", x"f902", x"f6d9", 
            x"f2e8", x"f0e5", x"f035", x"f293", 
            x"fa32", x"02a1", x"0481", x"fdee", 
            x"f149", x"e330", x"dd96", x"e774", 
            x"f847", x"0268", x"0396", x"033a", 
            x"085f", x"109f", x"1084", x"0426", 
            x"f426", x"e807", x"e28f", x"e54b", 
            x"eede", x"fa28", x"0147", x"01bb", 
            x"007f", x"0374", x"06e4", x"0470", 
            x"fed4", x"fed0", x"06b6", x"0e8a", 
            x"116c", x"11ea", x"0dff", x"04f5", 
            x"00e6", x"0542", x"0740", x"0217", 
            x"fdac", x"ff38", x"03d2", x"07b8", 
            x"09d0", x"0957", x"0623", x"03ac", 
            x"054e", x"07bd", x"074b", x"0712", 
            x"07f4", x"04ad", x"fdce", x"fc65", 
            x"03d5", x"0c99", x"0fa8", x"0cdb", 
            x"07d5", x"05f6", x"0937", x"0bcb", 
            x"08fd", x"0499", x"0499", x"0949", 
            x"0de0", x"1014", x"121b", x"1400", 
            x"13cd", x"1208", x"10c4", x"114f", 
            x"13fc", x"18cd", x"1be4", x"1598", 
            x"0794", x"fd83", x"fb85", x"fb04", 
            x"f7df", x"f641", x"fa4f", x"ff85", 
            x"ffb2", x"fe61", x"0255", x"085d", 
            x"087c", x"0354", x"000f", x"0071", 
            x"0055", x"fde2", x"fbc8", x"fcec", 
            x"02c0", x"0abd", x"0c92", x"0528", 
            x"fc94", x"fb5c", x"0242", x"0a9e", 
            x"0d1f", x"0815", x"fd45", x"f26f", 
            x"efc6", x"f3b0", x"f296", x"ea09", 
            x"e6f2", x"ef4d", x"f592", x"eed7", 
            x"e3dc", x"e02d", x"e34f", x"e916", 
            x"f019", x"f2b0", x"e95a", x"dc06", 
            x"dc62", x"e931", x"f0af", x"eefd", 
            x"ef8b", x"f54e", x"f842", x"f741", 
            x"fb97", x"0810", x"1247", x"123d", 
            x"0c01", x"0620", x"03e3", x"08c0", 
            x"1433", x"1cef", x"19fb", x"0fe1", 
            x"0ac4", x"0c25", x"0b69", x"0648", 
            x"059a", x"0fd6", x"1bab", x"1b26", 
            x"12ef", x"12b7", x"1934", x"182e", 
            x"0ebe", x"077d", x"0320", x"fb70", 
            x"f390", x"f240", x"f635", x"fb70", 
            x"014d", x"054c", x"00eb", x"f3ca", 
            x"e9df", x"ed17", x"f554", x"f407", 
            x"ead3", x"e7b0", x"ef51", x"f93e", 
            x"fd08", x"fb34", x"fc09", x"037e", 
            x"084e", x"01f3", x"f8ae", x"f6df", 
            x"f81d", x"f819", x"fc54", x"0274", 
            x"0078", x"fc81", x"055a", x"146c", 
            x"1920", x"16a6", x"16a6", x"1356", 
            x"07dc", x"fe0b", x"fd71", x"ffff", 
            x"fd08", x"f695", x"f5a1", x"f9b8", 
            x"f997", x"f3d2", x"ef90", x"f106", 
            x"f684", x"f928", x"f1bc", x"e5df", 
            x"e5c6", x"f2ab", x"f7ef", x"ea0f", 
            x"d9cc", x"db84", x"eb38", x"f6bc", 
            x"f9c9", x"fe9a", x"07ff", x"0f96", 
            x"1314", x"13c3", x"1088", x"0822", 
            x"0047", x"0287", x"0c63", x"0ff4", 
            x"08c4", x"ff55", x"faa2", x"fa39", 
            x"f9ec", x"f7d6", x"f725", x"f989", 
            x"fb3e", x"f9d8", x"f821", x"f6a2", 
            x"f1fc", x"ec4d", x"ec68", x"f17f", 
            x"f319", x"ef8f", x"ee6e", x"f1f5", 
            x"f398", x"f2f9", x"f87b", x"0194", 
            x"fee6", x"f117", x"ed1a", x"f932", 
            x"03a0", x"02dc", x"030c", x"0d3e", 
            x"197a", x"1bdd", x"12b8", x"0905", 
            x"0ad2", x"1579", x"1bf8", x"17ea", 
            x"0daa", x"04c2", x"00f4", x"032e", 
            x"0a7f", x"1091", x"112f", x"110e", 
            x"136e", x"150c", x"137d", x"0f43", 
            x"089d", x"026f", x"02da", x"08a0", 
            x"0a69", x"076d", x"05d5", x"045b", 
            x"0026", x"fd01", x"0019", x"070a", 
            x"0822", x"ffc2", x"f6fa", x"f970", 
            x"08e3", x"181f", x"14c2", x"ffab", 
            x"efd3", x"f29a", x"fad1", x"f9f9", 
            x"f6c0", x"fc99", x"0691", x"0b89", 
            x"0ece", x"142e", x"1663", x"1415", 
            x"120d", x"0e12", x"04ed", x"febb", 
            x"02a4", x"0a8e", x"0d58", x"09f8", 
            x"04de", x"0297", x"053b", x"08ad", 
            x"0264", x"f0e8", x"e667", x"f0f7", 
            x"01f7", x"0503", x"007c", x"03d4", 
            x"0a59", x"07cc", x"fdd4", x"f802"
        ),
        -- Block 12
        (
            x"fda4", x"0945", x"0ffc", x"0fd2", 
            x"0eab", x"0f9f", x"1052", x"0c67", 
            x"0400", x"fea4", x"ffdc", x"ffe6", 
            x"f802", x"ee1e", x"ece0", x"f5d2", 
            x"0082", x"05d5", x"066f", x"054b", 
            x"0267", x"fb0f", x"f0de", x"ec10", 
            x"ed66", x"eb49", x"e575", x"e780", 
            x"f41d", x"0026", x"0368", x"026c", 
            x"033f", x"0407", x"0198", x"fc03", 
            x"f4f8", x"f027", x"f1ee", x"f8d6", 
            x"fb3f", x"f45c", x"ed4b", x"ee93", 
            x"f2ec", x"f211", x"ec6e", x"e747", 
            x"e698", x"e857", x"e41f", x"d940", 
            x"d3fa", x"da70", x"e2fc", x"e472", 
            x"e250", x"e534", x"ef9c", x"fbfc", 
            x"0411", x"05e8", x"0242", x"fb88", 
            x"f530", x"f0fc", x"ef56", x"f098", 
            x"f455", x"fa83", x"0384", x"0e06", 
            x"1737", x"1d3a", x"20ab", x"20bf", 
            x"1910", x"0a69", x"fc69", x"f4c2", 
            x"f5dc", x"ff82", x"0b79", x"0fd8", 
            x"085f", x"fde8", x"fd4b", x"05d2", 
            x"0ba1", x"089e", x"00cd", x"f941", 
            x"f311", x"ef44", x"f201", x"fbb1", 
            x"025b", x"fd10", x"f291", x"f14b", 
            x"fa44", x"0108", x"0142", x"016f", 
            x"01c0", x"000b", x"02f3", x"0d14", 
            x"135b", x"0fe8", x"0e04", x"13ea", 
            x"13b3", x"0473", x"f47d", x"f10e", 
            x"f466", x"f7ea", x"ff53", x"0b2c", 
            x"12b9", x"1150", x"0da8", x"0d22", 
            x"0ca5", x"0c68", x"10ab", x"154a", 
            x"121c", x"0872", x"00a2", x"0010", 
            x"0695", x"0f7a", x"1421", x"13e9", 
            x"15f2", x"1d22", x"2063", x"1758", 
            x"0c08", x"0d3f", x"13d6", x"0f53", 
            x"020c", x"facd", x"fe19", x"0385", 
            x"04a5", x"0441", x"0382", x"fc9b", 
            x"f163", x"eede", x"f890", x"03a9", 
            x"0697", x"0076", x"f96e", x"faea", 
            x"0311", x"094a", x"08ca", x"03b3", 
            x"0261", x"06c6", x"06f3", x"fee3", 
            x"f7cc", x"f815", x"fb48", x"fa7a", 
            x"f5d3", x"f4f8", x"fdc8", x"0b2c", 
            x"0f3d", x"048a", x"f8a0", x"f931", 
            x"026b", x"0721", x"00bc", x"f6d7", 
            x"f522", x"f953", x"f7e0", x"f179", 
            x"f18b", x"f868", x"f9c0", x"f1c9", 
            x"ec69", x"f2ca", x"fc7a", x"fdd7", 
            x"fa7c", x"fa6f", x"fbe7", x"fc0e", 
            x"fbd6", x"f7af", x"ebf1", x"def0", 
            x"d872", x"d892", x"df0b", x"ebd1", 
            x"f755", x"f89c", x"f1a9", x"ed79", 
            x"f221", x"fa78", x"ff0e", x"fd16", 
            x"f45b", x"ea3d", x"eaab", x"f988", 
            x"08ea", x"0aaf", x"02c5", x"fd27", 
            x"fd44", x"ff61", x"01bc", x"05e7", 
            x"0931", x"04f8", x"f9cc", x"f02f", 
            x"ee54", x"f407", x"fbd1", x"feda", 
            x"fe49", x"01ad", x"0700", x"02f4", 
            x"f65d", x"f1bd", x"fba7", x"03f7", 
            x"fc45", x"ee64", x"eb80", x"f414", 
            x"fbf0", x"fcbe", x"fcb5", x"02c2", 
            x"0b42", x"0ebe", x"0ca1", x"098e", 
            x"0942", x"0d07", x"13fa", x"1882", 
            x"11e1", x"03d3", x"0071", x"0b88", 
            x"1341", x"0fc0", x"0ec8", x"1782", 
            x"1cfc", x"146e", x"07a7", x"059a", 
            x"0a73", x"084f", x"fe81", x"f513", 
            x"ed8d", x"e776", x"e6df", x"edc4", 
            x"f57b", x"f4d3", x"eea5", x"f024", 
            x"fa45", x"fe61", x"f865", x"f509", 
            x"f9f4", x"ff67", x"024a", x"0689", 
            x"099a", x"0643", x"026f", x"0799", 
            x"1052", x"0e74", x"030d", x"fe98", 
            x"0757", x"11fb", x"14e1", x"0fc0", 
            x"0386", x"f480", x"ed49", x"f16a", 
            x"f69a", x"f328", x"eb14", x"e8be", 
            x"eda4", x"f2c0", x"f549", x"f7bb", 
            x"f920", x"f706", x"f53a", x"f940", 
            x"0092", x"04cc", x"0548", x"0640", 
            x"0b09", x"1182", x"12b5", x"107b", 
            x"1763", x"260e", x"2a68", x"204d", 
            x"1784", x"173e", x"16d7", x"1203", 
            x"0fae", x"15f2", x"1e5d", x"1e12", 
            x"1791", x"12a3", x"0d2f", x"0591", 
            x"009d", x"ff3b", x"fcbd", x"f79c", 
            x"f4b1", x"f9b5", x"0449", x"0832", 
            x"ffc0", x"f6fa", x"f81b", x"fb32", 
            x"f7d9", x"f3da", x"f7db", x"036b", 
            x"0f51", x"1437", x"10f3", x"0c98", 
            x"0d30", x"108f", x"1090", x"0a56", 
            x"0327", x"0331", x"07db", x"07e5", 
            x"0446", x"0555", x"0b98", x"0f2f", 
            x"0c7c", x"075d", x"063c", x"0c05", 
            x"126b", x"0f99", x"05d2", x"0082", 
            x"025f", x"05f2", x"090c", x"0b54", 
            x"0890", x"ffc2", x"f99f", x"fad6", 
            x"fdd5", x"0235", x"0a60", x"0de1", 
            x"051f", x"f9fe", x"fa6d", x"02b3", 
            x"0571", x"02e3", x"03d2", x"066e", 
            x"06aa", x"092e", x"0de1", x"0bb1", 
            x"01b5", x"f9ea", x"f844", x"f666", 
            x"f378", x"f396", x"f263", x"ed8a", 
            x"ee5a", x"f86e", x"0110", x"ffcc", 
            x"fb70", x"fe93", x"0572", x"0485", 
            x"fe12", x"fe9e", x"0644", x"0a08", 
            x"07a4", x"0418", x"ff33", x"f78e", 
            x"f15b", x"f08c", x"f339", x"f50e", 
            x"f553", x"f762", x"faa5", x"f9a3", 
            x"f5df", x"f79a", x"fe85", x"00bd", 
            x"f949", x"ed07", x"e4dd", x"e723", 
            x"f1a1", x"f99b", x"f8af", x"f529", 
            x"f5ef", x"f8f0", x"fb05", x"fdd4", 
            x"021a", x"0583", x"06f3", x"08dc", 
            x"0e4f", x"175e", x"2209", x"27f2", 
            x"224b", x"174a", x"15c0", x"1ed6", 
            x"21a0", x"15cf", x"084f", x"044a", 
            x"0640", x"07a2", x"056e", x"fcf1", 
            x"efe8", x"e761", x"e79a", x"e8bb", 
            x"e3f4", x"df97", x"e5f0", x"f3f7", 
            x"fcf7", x"fca0", x"f7c8", x"f276", 
            x"f018", x"f499", x"fc6b", x"ffc3", 
            x"fe85", x"fbc8", x"f82e", x"f5b5", 
            x"f46d", x"f206", x"f19d", x"f7b7", 
            x"ff33", x"ffc7", x"fc5f", x"fe92", 
            x"0839", x"11f3", x"133f", x"09dd", 
            x"fb3d", x"efa4", x"ec8c", x"f0b9", 
            x"f4c8", x"f339", x"eed4", x"ef73", 
            x"f7d5", x"ffbb", x"ff80", x"fbc5", 
            x"fd43", x"029f", x"03f7", x"0043", 
            x"fd83", x"fedb", x"ff24", x"f812", 
            x"f2e6", x"00ff", x"1ada", x"23be", 
            x"1586", x"06b7", x"0670", x"0e48", 
            x"1554", x"1c7c", x"205b", x"17ec", 
            x"0a5f", x"0879", x"0fb7", x"0f72", 
            x"0438", x"fb80", x"fef9", x"0638", 
            x"033a", x"f70f", x"ee45", x"ef36", 
            x"f5ff", x"fbbe", x"f9b4", x"edf9", 
            x"e397", x"e888", x"f8d6", x"0198", 
            x"f9fd", x"ec8f", x"e7f9", x"ef89", 
            x"f88d", x"f5fc", x"ea74", x"e5e5", 
            x"ef24", x"fbba", x"0052", x"0027", 
            x"042b", x"09a4", x"063a", x"fb33", 
            x"f575", x"fa13", x"ff62", x"fd87", 
            x"f9c5", x"f960", x"f956", x"f9e0", 
            x"ff3c", x"0431", x"0251", x"01ae", 
            x"0b28", x"14f6", x"116d", x"0568", 
            x"ffc3", x"04d7", x"0a9f", x"06db", 
            x"fc59", x"f581", x"f5c2", x"f828", 
            x"f9bf", x"fc41", x"fe37", x"faa5", 
            x"f2eb", x"f0c2", x"f7ae", x"fad9", 
            x"efaf", x"e275", x"e4c4", x"f088", 
            x"f288", x"e9b9", x"e42f", x"e4c7", 
            x"e4af", x"e8e9", x"f832", x"0595", 
            x"01c8", x"f40d", x"ede1", x"f2eb", 
            x"f85d", x"f755", x"f4f6", x"f43c", 
            x"f219", x"f159", x"f790", x"03df", 
            x"10ba", x"1764", x"1493", x"0c0a", 
            x"044d", x"021f", x"0531", x"07f2", 
            x"0482", x"fa0c", x"f00f", x"eeff", 
            x"f499", x"fbb0", x"0602", x"0f95", 
            x"0c11", x"fb58", x"ec47", x"e6f4", 
            x"e640", x"e5fe", x"e922", x"f264", 
            x"feab", x"07c6", x"0a33", x"088e", 
            x"082b", x"0a1a", x"0a40", x"06ba", 
            x"035d", x"03df", x"06c6", x"08ae", 
            x"0a8b", x"0f34", x"1550", x"1a97", 
            x"1ede", x"1f33", x"19d3", x"1502", 
            x"16cc", x"1c6d", x"1ed3", x"1b18", 
            x"13c7", x"0ab7", x"0102", x"ff6f", 
            x"0c0f", x"177d", x"0d9f", x"f4ec", 
            x"e773", x"f020", x"fda4", x"fcfa", 
            x"f383", x"f1ca", x"f8c5", x"fda4", 
            x"fe60", x"ffa2", x"fef5", x"fa11", 
            x"f986", x"03c7", x"1137", x"1625", 
            x"1069", x"09e6", x"0f05", x"1e42", 
            x"2802", x"2508", x"1f33", x"2080", 
            x"274f", x"2b84", x"273a", x"1b8e", 
            x"0f19", x"08d8", x"0aa9", x"1117", 
            x"186c", x"1b10", x"12d9", x"0402", 
            x"fbea", x"00d2", x"08c2", x"0560", 
            x"f6ec", x"ecc9", x"f17c", x"fab7", 
            x"fa37", x"f537", x"f7a5", x"fc3a", 
            x"f6df", x"ec4f", x"ed3b", x"fd2c", 
            x"0ae7", x"0944", x"018e", x"007a", 
            x"0517", x"096e", x"0970", x"03b7", 
            x"fc95", x"fdde", x"0b79", x"188f", 
            x"161a", x"0938", x"016d", x"0297", 
            x"07cf", x"0d32", x"0fea", x"0ec7", 
            x"0cc1", x"0c2d", x"08c5", x"ff85", 
            x"f5cc", x"f1a0", x"f1a8", x"f178", 
            x"f099", x"f086", x"ef26", x"ec80", 
            x"ee2d", x"f430", x"f700", x"f3ac", 
            x"ef7b", x"ed08", x"e88b", x"e2bf", 
            x"e448", x"f0d8", x"fcf1", x"fba9", 
            x"f392", x"f5f4", x"0396", x"0b93", 
            x"0560", x"feac", x"05ad", x"0eb4", 
            x"0629", x"f430", x"f113", x"fef3", 
            x"0af4", x"0a3c", x"0097", x"f5aa", 
            x"efe9", x"f107", x"f397", x"f318", 
            x"f2b1", x"f4c7", x"f47a", x"effa", 
            x"eef8", x"f4fa", x"f7cd", x"ef8d", 
            x"e4b3", x"e312", x"ea95", x"f389", 
            x"f7e0", x"f7c3", x"f728", x"f513", 
            x"ef99", x"ed04", x"f093", x"efdd", 
            x"e4d6", x"db5d", x"e072", x"efe3", 
            x"fab5", x"fa21", x"f4e4", x"f55c", 
            x"00fa", x"1229", x"1a09", x"1337", 
            x"0b38", x"0ee9", x"1646", x"0ed9", 
            x"f9d4", x"ee02", x"f537", x"feea", 
            x"fc4e", x"f34d", x"ee26", x"eeb1", 
            x"f55e", x"0195", x"0a0e", x"0530", 
            x"f800", x"f11e", x"f7e8", x"04fa", 
            x"0943", x"002c", x"f612", x"f414", 
            x"f543", x"f44e", x"f335", x"f59b", 
            x"fa87", x"fbc0", x"f750", x"f449", 
            x"f58d", x"f2f0", x"eb1b", x"ec6f", 
            x"fceb", x"0b3a", x"071c", x"f75a", 
            x"ef8f", x"fa38", x"0cae", x"13ad", 
            x"0c88", x"04bc", x"045e", x"0843", 
            x"09f1", x"052d", x"fcd6", x"fac3", 
            x"042c", x"10ec", x"1339", x"0808", 
            x"fc88", x"fc46", x"0138", x"013d", 
            x"fdb8", x"fa27", x"f2fe", x"e986", 
            x"e990", x"f6bd", x"048e", x"08c9", 
            x"0711", x"0a0b", x"120c", x"1268", 
            x"08b5", x"0317", x"0780", x"0c8f", 
            x"0b9c", x"06dc", x"0350", x"013e", 
            x"fced", x"f9e3", x"fd7a", x"010e", 
            x"ff26", x"fe93", x"0060", x"fddc", 
            x"fb59", x"ff78", x"02e0", x"fdad", 
            x"f606", x"f620", x"fcda", x"0266", 
            x"0601", x"0a99", x"0d56", x"0b9e", 
            x"092d", x"0628", x"fe47", x"f580", 
            x"f3f7", x"fa13", x"03b3", x"0cd7", 
            x"12d0", x"166d", x"179b", x"1436", 
            x"0f17", x"0d62", x"0ea5", x"106a", 
            x"1518", x"1c13", x"1e21", x"1b03", 
            x"19b3", x"1baa", x"1c43", x"171e", 
            x"0eb6", x"0a38", x"08ad", x"05c4", 
            x"0531", x"0978", x"0d2d", x"0d09", 
            x"0cd6", x"0ede", x"0efb", x"0a68", 
            x"03df", x"fd9c", x"f7a9", x"f211", 
            x"f022", x"f63e", x"0061", x"0456", 
            x"0107", x"ff55", x"01e0", x"ff8b", 
            x"f581", x"f278", x"00cf", x"1277", 
            x"1344", x"057a", x"fe32", x"0722", 
            x"1278", x"1211", x"0a6f", x"08ff", 
            x"116e", x"19a1", x"1830", x"12ce", 
            x"13f3", x"1a3d", x"1ee7", x"200b", 
            x"2060", x"2395", x"2689", x"20db", 
            x"1510", x"1015", x"1612", x"1d15", 
            x"1c24", x"14ad", x"0c5d", x"07ac", 
            x"0863", x"0917", x"023b", x"f8f0", 
            x"f79b", x"fa41", x"f6ab", x"ee7e"
        ),
        -- Block 11
        (
            x"eaf2", x"edea", x"ef24", x"eb45", 
            x"e87e", x"e60a", x"df28", x"da25", 
            x"dcef", x"e4f8", x"f0ac", x"fb34", 
            x"f775", x"e494", x"d963", x"e5f1", 
            x"f998", x"fb7b", x"ef79", x"eb7e", 
            x"f246", x"f0ce", x"e131", x"d80d", 
            x"e2dc", x"f370", x"f769", x"eff0", 
            x"ec06", x"f375", x"fce4", x"fd0a", 
            x"f783", x"f698", x"fc76", x"023f", 
            x"02a3", x"fcac", x"f206", x"eb7e", 
            x"f112", x"fbd0", x"fcb3", x"f205", 
            x"eadb", x"eee2", x"f370", x"f48f", 
            x"fac3", x"0486", x"0947", x"08bc", 
            x"062a", x"032e", x"0279", x"06d8", 
            x"0ea0", x"111e", x"0a2a", x"0341", 
            x"01e3", x"fd8b", x"f5b4", x"f99a", 
            x"092b", x"0aec", x"f569", x"e5b8", 
            x"f2b9", x"0a85", x"10dc", x"0413", 
            x"f692", x"f359", x"f84a", x"0044", 
            x"0520", x"00f7", x"f8a7", x"f9c7", 
            x"04d4", x"09a8", x"0200", x"f9ce", 
            x"f888", x"f8b2", x"f79f", x"f8cb", 
            x"fbc9", x"fea5", x"02f9", x"0820", 
            x"09f7", x"096f", x"0b82", x"0d5a", 
            x"07fc", x"ffd6", x"ff50", x"0281", 
            x"fc57", x"f078", x"efcb", x"fa5d", 
            x"ffce", x"fd24", x"fdd8", x"ffc6", 
            x"f734", x"ebea", x"ed26", x"f4a5", 
            x"f2cb", x"e8f4", x"e690", x"f1a0", 
            x"feef", x"0590", x"0917", x"0a17", 
            x"03b6", x"f9d1", x"f62a", x"fc96", 
            x"080a", x"1005", x"12de", x"1426", 
            x"15c9", x"18cd", x"18ec", x"1098", 
            x"06b6", x"06ab", x"0be1", x"08ce", 
            x"ff53", x"fd4b", x"03e9", x"0854", 
            x"0781", x"0634", x"0486", x"ff5a", 
            x"f95b", x"f5de", x"f2ab", x"edb8", 
            x"e6c4", x"df7c", x"de9f", x"e7e4", 
            x"f23a", x"f233", x"e7f4", x"dfe0", 
            x"e6b3", x"f644", x"fc36", x"f79e", 
            x"f68e", x"fdd5", x"0a62", x"1783", 
            x"1bef", x"15ac", x"11bc", x"179e", 
            x"1dcf", x"1999", x"0c14", x"0121", 
            x"03ff", x"1231", x"1dec", x"1c47", 
            x"0cf3", x"faef", x"f315", x"f690", 
            x"fad5", x"f981", x"fa95", x"003c", 
            x"fd8a", x"f28d", x"ef75", x"f5f5", 
            x"f81e", x"f247", x"f035", x"fa4f", 
            x"08f1", x"0d94", x"05e9", x"fee3", 
            x"01d8", x"05e6", x"0027", x"f845", 
            x"fae2", x"01d3", x"0172", x"ff59", 
            x"0334", x"0810", x"0914", x"07e2", 
            x"0428", x"fc8d", x"f417", x"f0b5", 
            x"f537", x"fb0d", x"f843", x"ef0a", 
            x"ee46", x"fcde", x"0ba8", x"07e0", 
            x"f82f", x"f197", x"f793", x"fe45", 
            x"ff6e", x"fd5b", x"f979", x"f629", 
            x"fbcf", x"0cec", x"1c90", x"1b8c", 
            x"0a77", x"fba1", x"fe30", x"08cd", 
            x"05d2", x"f480", x"ed8e", x"fdec", 
            x"1247", x"144d", x"083e", x"0137", 
            x"0460", x"06b5", x"001e", x"f3fb", 
            x"e8fd", x"e2be", x"e4c6", x"eef1", 
            x"fa3c", x"0061", x"0168", x"0091", 
            x"fe67", x"fafb", x"f958", x"f779", 
            x"f05a", x"eb12", x"f2f4", x"017d", 
            x"0776", x"0641", x"0a78", x"13b4", 
            x"1483", x"0c58", x"0a7e", x"1269", 
            x"1724", x"132c", x"0d80", x"0ac4", 
            x"08b1", x"0936", x"11da", x"1e1a", 
            x"20b1", x"14d3", x"07c3", x"09ee", 
            x"1b62", x"295b", x"218b", x"09d6", 
            x"fa79", x"fc8a", x"0146", x"fecc", 
            x"fd39", x"0234", x"05c3", x"011f", 
            x"f928", x"f732", x"fca4", x"02a0", 
            x"0425", x"0311", x"0385", x"0587", 
            x"05d3", x"0494", x"0613", x"0a85", 
            x"0bb9", x"0628", x"fe7a", x"f9ed", 
            x"f7b6", x"f87f", x"fe34", x"048e", 
            x"0752", x"0750", x"0571", x"01f5", 
            x"000c", x"021b", x"04f3", x"01a6", 
            x"f52a", x"e868", x"e6e8", x"f051", 
            x"fc3e", x"01d3", x"fcdd", x"f61c", 
            x"fbdd", x"0ae2", x"10cb", x"06f1", 
            x"f9e9", x"f653", x"fb9f", x"02b4", 
            x"05df", x"0020", x"f4f1", x"f34d", 
            x"fdda", x"0496", x"0044", x"faf4", 
            x"fda3", x"0517", x"095a", x"098e", 
            x"0a04", x"0a39", x"04cd", x"f882", 
            x"ec45", x"e710", x"e7d3", x"e977", 
            x"ea87", x"ee22", x"f6a9", x"fef0", 
            x"ff9f", x"fbdc", x"fbf1", x"fd6c", 
            x"fc5d", x"fedc", x"06ef", x"0c65", 
            x"0a00", x"0495", x"03ed", x"08db", 
            x"0ec4", x"1525", x"19b9", x"1521", 
            x"0a75", x"06ff", x"0f4d", x"178f", 
            x"12e9", x"0421", x"f7f7", x"f605", 
            x"fb56", x"0113", x"04c3", x"068a", 
            x"0345", x"fac0", x"f6b7", x"fb28", 
            x"fecc", x"ff7c", x"0530", x"0e73", 
            x"120c", x"0c93", x"06a9", x"0b03", 
            x"127b", x"0ec8", x"021b", x"f934", 
            x"f94e", x"fc92", x"fdf4", x"0171", 
            x"09aa", x"1121", x"117c", x"0a89", 
            x"ff57", x"f29a", x"ec2a", x"f4b2", 
            x"04d1", x"0a93", x"0345", x"fe13", 
            x"04a0", x"0e6c", x"0f28", x"06f8", 
            x"fe20", x"fb26", x"fda3", x"fe97", 
            x"fb04", x"f7fb", x"f6e6", x"f5a4", 
            x"f51c", x"f394", x"ee59", x"ea6d", 
            x"edd5", x"f679", x"fda9", x"fe4f", 
            x"fd29", x"02da", x"0841", x"ff54", 
            x"ec0e", x"e03b", x"e53e", x"f1cb", 
            x"f788", x"f657", x"f63e", x"f5e4", 
            x"f29c", x"f1ef", x"f69a", x"fa36", 
            x"f542", x"ea69", x"e747", x"f24f", 
            x"ffe7", x"057e", x"04cd", x"0245", 
            x"ff9a", x"fdc2", x"fc7e", x"f905", 
            x"f440", x"f4fa", x"fb17", x"fe21", 
            x"fb53", x"f628", x"f19f", x"eecf", 
            x"ee3d", x"f020", x"f138", x"ebc0", 
            x"e2a2", x"deee", x"e0ef", x"e5fc", 
            x"f23d", x"0213", x"0549", x"f6dc", 
            x"e872", x"eaca", x"f536", x"f74e", 
            x"f59a", x"fb5a", x"00ac", x"facc", 
            x"f2bd", x"f669", x"0273", x"08da", 
            x"05b7", x"0296", x"0956", x"1731", 
            x"1e59", x"1612", x"06b9", x"fe2a", 
            x"fcdb", x"fbea", x"fc44", x"fea4", 
            x"fa39", x"ebd9", x"e308", x"ef05", 
            x"00ef", x"010c", x"f784", x"f689", 
            x"faf5", x"0059", x"084f", x"09e0", 
            x"ffcd", x"f691", x"f853", x"ff15", 
            x"04f8", x"0cab", x"10e9", x"0877", 
            x"fcde", x"fe24", x"07a6", x"0c17", 
            x"0be5", x"0d6c", x"0f76", x"1038", 
            x"1160", x"1115", x"0d7f", x"09d4", 
            x"080c", x"06de", x"066f", x"06e8", 
            x"07a7", x"071e", x"0359", x"ffd7", 
            x"fddf", x"f436", x"e43a", x"e0a3", 
            x"eadd", x"ed84", x"e288", x"d95e", 
            x"dca0", x"eabd", x"fc26", x"070e", 
            x"05fc", x"fd3d", x"f9ca", x"01b2", 
            x"0a98", x"0952", x"0101", x"ff96", 
            x"09ee", x"1373", x"1297", x"0ecc", 
            x"14af", x"251e", x"31c6", x"2d3f", 
            x"1d6c", x"16d2", x"1f61", x"2632", 
            x"2066", x"177e", x"156b", x"17ad", 
            x"1843", x"150a", x"0fb3", x"0b99", 
            x"0837", x"008d", x"f2ea", x"e71f", 
            x"e826", x"f1c5", x"f477", x"ef9e", 
            x"ee06", x"efde", x"ee41", x"ea43", 
            x"eac3", x"ee0b", x"eca0", x"e8ba", 
            x"e9d1", x"efaa", x"f550", x"f706", 
            x"f341", x"f0b5", x"faf6", x"1226", 
            x"28b5", x"3181", x"2bd7", x"2209", 
            x"1c38", x"1c3b", x"20b0", x"208e", 
            x"1649", x"0b54", x"0807", x"0989", 
            x"0ba5", x"0cf7", x"0dec", x"0e6b", 
            x"0b72", x"07db", x"0aba", x"10dc", 
            x"12c9", x"0f73", x"05c9", x"f99c", 
            x"f544", x"fae7", x"026c", x"025e", 
            x"f7e8", x"ea1e", x"e26c", x"e342", 
            x"e9d2", x"f311", x"fd25", x"0740", 
            x"0d9c", x"0c72", x"0944", x"0ad2", 
            x"0b62", x"030c", x"f5f3", x"ebde", 
            x"e90c", x"f119", x"ffa6", x"08a8", 
            x"0760", x"04e1", x"0b2d", x"1444", 
            x"151d", x"0d66", x"02c0", x"fbec", 
            x"fddf", x"05ac", x"0b2f", x"0a3a", 
            x"04f3", x"020c", x"0372", x"0204", 
            x"fce0", x"fbeb", x"0185", x"06ad", 
            x"0499", x"fda9", x"f957", x"fd37", 
            x"0673", x"0acd", x"0782", x"04e0", 
            x"073f", x"0c66", x"11f5", x"14c1", 
            x"1189", x"08da", x"01b9", x"027f", 
            x"0726", x"07ab", x"042d", x"018f", 
            x"004d", x"ff61", x"024c", x"08de", 
            x"0a98", x"03ef", x"fbc8", x"f797", 
            x"f4b9", x"eff1", x"ecb9", x"ef89", 
            x"f336", x"ef58", x"eaaf", x"f2f3", 
            x"0387", x"0ac7", x"018c", x"f286", 
            x"ecae", x"f2b4", x"fe9b", x"0a7d", 
            x"0bb3", x"fea1", x"f6c0", x"0145", 
            x"0b39", x"04e7", x"fe44", x"065f", 
            x"143f", x"1d05", x"1fd8", x"1ead", 
            x"1dd4", x"1f8d", x"1e8b", x"1b48", 
            x"1c8a", x"217a", x"246c", x"1bd3", 
            x"034a", x"ee09", x"f10c", x"016b", 
            x"0834", x"039a", x"fe84", x"fd4e", 
            x"fdf7", x"fd6a", x"fa0b", x"f71a", 
            x"f432", x"e9b0", x"db6c", x"d6c3", 
            x"da0c", x"da9a", x"dbb9", x"e46b", 
            x"ecd1", x"e88c", x"db4c", x"d744", 
            x"e5ab", x"f7d8", x"fbae", x"f651", 
            x"f5cd", x"fa2d", x"fe70", x"02c2", 
            x"05e4", x"0490", x"0046", x"fc88", 
            x"f7a8", x"f07c", x"eb5c", x"ee1d", 
            x"fa3b", x"03cb", x"fe35", x"f159", 
            x"eb24", x"ee3e", x"f6b4", x"fbc4", 
            x"f5dc", x"e80c", x"dc7d", x"db24", 
            x"e1b6", x"e5d2", x"e1c6", x"d9f3", 
            x"d538", x"d18c", x"c9f3", x"c589", 
            x"d0bf", x"e860", x"f70e", x"ef81", 
            x"de90", x"dc03", x"ee21", x"ff96", 
            x"fc0c", x"ed3f", x"e864", x"ec83", 
            x"ed9f", x"ee41", x"f499", x"fe6e", 
            x"0672", x"0514", x"f716", x"e9a1", 
            x"eb8f", x"f72d", x"fd27", x"fc11", 
            x"000f", x"0c79", x"111b", x"04ea", 
            x"f958", x"f9b1", x"f8a2", x"f027", 
            x"ed86", x"f681", x"00bc", x"05cf", 
            x"082c", x"0812", x"0620", x"06c9", 
            x"0b56", x"0eaa", x"09ee", x"000c", 
            x"fe95", x"0a57", x"1b52", x"2718", 
            x"2496", x"1956", x"14bd", x"1441", 
            x"0d4a", x"06e7", x"0cc0", x"1935", 
            x"1ce2", x"1354", x"07be", x"0595", 
            x"0a21", x"0b7c", x"091d", x"097b", 
            x"0808", x"faef", x"eb71", x"ec4b", 
            x"fc7b", x"0a5a", x"0d67", x"0e86", 
            x"12d3", x"1432", x"14ac", x"1b29", 
            x"2203", x"1ec8", x"1172", x"04ee", 
            x"02f2", x"077d", x"07f9", x"056b", 
            x"0640", x"089c", x"0c8c", x"132f", 
            x"11a2", x"013c", x"ef50", x"e9be", 
            x"ee56", x"f487", x"fb88", x"0301", 
            x"0306", x"fd37", x"00ed", x"0f4d", 
            x"1420", x"0721", x"fad8", x"0111", 
            x"13fd", x"211c", x"2129", x"1f4b", 
            x"25c9", x"2ad7", x"23db", x"18df", 
            x"13db", x"1772", x"1ea5", x"1d1b", 
            x"12f4", x"105c", x"18ef", x"1c03", 
            x"129c", x"08dd", x"02e2", x"fc45", 
            x"f7ab", x"f4d7", x"ed05", x"e2b8", 
            x"de97", x"e1f1", x"e8cf", x"ed40", 
            x"eade", x"e777", x"e5cf", x"de20", 
            x"d8a4", x"e4d9", x"f484", x"ef73", 
            x"dffb", x"e53b", x"01e2", x"17e3", 
            x"1645", x"0c44", x"09a6", x"0a33", 
            x"085a", x"09b9", x"0eef", x"1241", 
            x"1567", x"19e1", x"1c26", x"1b54", 
            x"177c", x"0f50", x"05fa", x"0416", 
            x"0af2", x"0c38", x"ff74", x"f319", 
            x"f5eb", x"00ea", x"0400", x"fd23", 
            x"f679", x"f298", x"f23e", x"fc91", 
            x"0c9c", x"11a9", x"08af", x"fd98", 
            x"f7d3", x"f7a1", x"fbc3", x"fba1", 
            x"eedd", x"e0ed", x"e565", x"f983", 
            x"090b", x"0938", x"01c0", x"fde8", 
            x"fd80", x"fcc4", x"fd0f", x"01eb", 
            x"0b40", x"12d5", x"120d", x"0c45", 
            x"0bfb", x"1399", x"1897", x"14cd", 
            x"0ff1", x"1189", x"180e", x"1fc0", 
            x"22c7", x"1993", x"0849", x"fd80", 
            x"0023", x"0808", x"0791", x"fce0"
        ),
        -- Block 10
        (
            x"f456", x"f859", x"05c4", x"0dd1", 
            x"067e", x"f845", x"f28f", x"fa6e", 
            x"04b5", x"033f", x"fc16", x"fadc", 
            x"f9be", x"f1e8", x"e985", x"e8c9", 
            x"ef6f", x"f684", x"f99d", x"fa11", 
            x"fa94", x"fae0", x"fa8b", x"fd47", 
            x"039c", x"055d", x"0005", x"0024", 
            x"0b04", x"1367", x"1062", x"0952", 
            x"0812", x"0c4d", x"0f1b", x"0ba8", 
            x"05cd", x"04cb", x"08a0", x"0bb7", 
            x"0bc2", x"0c77", x"0c55", x"05a4", 
            x"fd05", x"f89d", x"f866", x"fe2c", 
            x"0627", x"0403", x"f86d", x"f136", 
            x"f308", x"f7c9", x"fa2f", x"fa1a", 
            x"f89c", x"f762", x"f8ad", x"fb7c", 
            x"fdbd", x"fe28", x"fc8a", x"fc75", 
            x"0066", x"02a4", x"fc1f", x"f403", 
            x"f766", x"02f9", x"09fe", x"0abe", 
            x"0bce", x"0f29", x"12ab", x"13c0", 
            x"1121", x"0ec4", x"0f6e", x"0dc4", 
            x"0462", x"f6fb", x"eedf", x"ee38", 
            x"edc2", x"eba5", x"ee81", x"f34b", 
            x"eee2", x"e56d", x"e6ab", x"f2c3", 
            x"fac3", x"f675", x"eb69", x"e136", 
            x"d810", x"d2d1", x"d9ac", x"e7b7", 
            x"ef4b", x"ee37", x"e8f8", x"e50c", 
            x"e8c5", x"f39c", x"0047", x"072c", 
            x"008f", x"f780", x"0032", x"11aa", 
            x"14d2", x"0b84", x"07ad", x"0c88", 
            x"0a46", x"fe8f", x"fd1a", x"06c5", 
            x"0669", x"fc64", x"ff24", x"1074", 
            x"13b0", x"fc06", x"e328", x"dee6", 
            x"e377", x"e0e0", x"ddcb", x"e17c", 
            x"e51b", x"e683", x"ea74", x"eee1", 
            x"edbc", x"e971", x"eb69", x"f1aa", 
            x"f01d", x"e9ef", x"e9f7", x"ec7c", 
            x"ef1d", x"f741", x"0003", x"ff21", 
            x"f4a4", x"ec10", x"f4d3", x"0e37", 
            x"2123", x"1d47", x"0ee7", x"0aa7", 
            x"0e2d", x"0cb4", x"091e", x"0aa8", 
            x"0c82", x"06ca", x"fce1", x"f9ee", 
            x"00f3", x"0b13", x"13c2", x"182f", 
            x"1223", x"043a", x"027e", x"13e5", 
            x"1e61", x"1056", x"fa83", x"f1d3", 
            x"f6d3", x"006c", x"09f0", x"0e58", 
            x"08d9", x"ff28", x"fc31", x"012f", 
            x"02bb", x"fc1d", x"fa14", x"ff98", 
            x"0033", x"fc08", x"fe17", x"0430", 
            x"02a2", x"fc61", x"fe33", x"0720", 
            x"0be1", x"066b", x"fae7", x"f4c9", 
            x"f9b6", x"0168", x"02bf", x"ffd9", 
            x"fea1", x"fcbb", x"f55a", x"f0f8", 
            x"fac8", x"0bc9", x"12fe", x"0b4c", 
            x"fcd2", x"f231", x"f323", x"fb54", 
            x"fe0d", x"f7ce", x"ed6b", x"e4e7", 
            x"e526", x"f1e3", x"0383", x"0cd9", 
            x"0bca", x"08fd", x"0aa7", x"10ec", 
            x"1821", x"1ab2", x"1786", x"10e6", 
            x"0764", x"0078", x"0437", x"0c1c", 
            x"083b", x"f854", x"ef7b", x"f918", 
            x"0759", x"0885", x"ffae", x"f7fc", 
            x"f2f0", x"f149", x"f57b", x"fa2f", 
            x"f76c", x"ef2b", x"eda4", x"f781", 
            x"007c", x"01b5", x"036b", x"05b1", 
            x"ff73", x"f540", x"f45c", x"fc91", 
            x"00a4", x"f889", x"edd5", x"ec12", 
            x"f0b3", x"f8ec", x"0232", x"ff29", 
            x"f169", x"ed7b", x"f315", x"f2a1", 
            x"ee57", x"f22e", x"fcb4", x"0496", 
            x"0893", x"0af5", x"07af", x"fe17", 
            x"f698", x"f1c4", x"ea7e", x"e639", 
            x"ec89", x"fc4d", x"0d2f", x"1371", 
            x"0c16", x"ffba", x"f634", x"f4ec", 
            x"fb08", x"fc71", x"f5c5", x"f4ed", 
            x"ff03", x"0b57", x"15df", x"1d39", 
            x"1b68", x"0f83", x"0260", x"fbb9", 
            x"fd1e", x"0462", x"0a6c", x"0ae7", 
            x"0e16", x"1784", x"1b79", x"16f6", 
            x"17c5", x"2015", x"1e78", x"0f32", 
            x"0878", x"1137", x"11c4", x"03e8", 
            x"fe46", x"06f4", x"0ccf", x"0610", 
            x"fad6", x"f908", x"ff59", x"003b", 
            x"fc34", x"f97c", x"f311", x"eaee", 
            x"ebf7", x"f5b8", x"fdcf", x"fce0", 
            x"f83f", x"faae", x"00eb", x"01a2", 
            x"0060", x"0686", x"1198", x"143a", 
            x"09e3", x"0165", x"08b9", x"15dd", 
            x"1734", x"0e34", x"0708", x"075d", 
            x"1079", x"1fa4", x"260c", x"1bf0", 
            x"12e8", x"1960", x"250a", x"27e9", 
            x"1fba", x"12ef", x"0942", x"028d", 
            x"fedd", x"01e2", x"063d", x"00d5", 
            x"f224", x"ea2e", x"f60b", x"09f5", 
            x"0fc5", x"0629", x"fcdb", x"fcd9", 
            x"056b", x"0fbc", x"0d23", x"f888", 
            x"e687", x"ef67", x"0a49", x"12b9", 
            x"fcea", x"e949", x"f00e", x"fe7c", 
            x"fdb2", x"f8d9", x"0232", x"0e1a", 
            x"0a0a", x"fdf5", x"f991", x"fde6", 
            x"0244", x"007c", x"fcd0", x"fe4a", 
            x"027d", x"04a6", x"06be", x"0860", 
            x"0554", x"ff59", x"fc82", x"fe44", 
            x"0019", x"03be", x"0d38", x"14c3", 
            x"1245", x"0ea6", x"1687", x"20bf", 
            x"198f", x"06b0", x"0411", x"1587", 
            x"1f9b", x"1408", x"0165", x"f5b7", 
            x"f5a9", x"0295", x"12be", x"176d", 
            x"0da2", x"ffed", x"fa3d", x"fd1c", 
            x"ff23", x"fcf2", x"fbda", x"fbad", 
            x"f911", x"f94a", x"fdad", x"fd2c", 
            x"f4fa", x"ea8a", x"e265", x"e365", 
            x"f0c0", x"fe6f", x"ffbd", x"f867", 
            x"f1a6", x"f083", x"f83c", x"ffbd", 
            x"f64c", x"e251", x"df88", x"f095", 
            x"f595", x"e6a8", x"e48c", x"f965", 
            x"0833", x"040e", x"feb1", x"026c", 
            x"065c", x"043e", x"0225", x"0456", 
            x"0625", x"055a", x"0708", x"0c43", 
            x"0dbd", x"09fe", x"06c7", x"091c", 
            x"14ee", x"221c", x"1f22", x"0fc2", 
            x"09a5", x"0f3a", x"0fb3", x"075f", 
            x"0167", x"fdc0", x"f8a8", x"f9ff", 
            x"ff37", x"f8f4", x"ee2a", x"f474", 
            x"02a1", x"fcb1", x"e58e", x"db6a", 
            x"e3cf", x"e5c7", x"dc05", x"da61", 
            x"e3b0", x"e896", x"e6f8", x"e6c2", 
            x"e576", x"de7d", x"da57", x"dde3", 
            x"df55", x"debc", x"e908", x"fbaa", 
            x"0415", x"ff3a", x"fce0", x"030b", 
            x"0898", x"070e", x"ff24", x"f3ad", 
            x"e9b9", x"e603", x"ea1e", x"f3d9", 
            x"fbed", x"fc00", x"f696", x"f2b6", 
            x"f24e", x"f3ea", x"f8fa", x"0131", 
            x"0870", x"0c1c", x"0f15", x"13fe", 
            x"1678", x"1373", x"0e4f", x"0859", 
            x"026b", x"feed", x"fe55", x"0677", 
            x"1762", x"22b7", x"1e79", x"0c22", 
            x"fc7e", x"03e5", x"1615", x"15b7", 
            x"05bb", x"ff8c", x"040d", x"0226", 
            x"0078", x"0fbf", x"224f", x"203c", 
            x"10a6", x"0a50", x"106b", x"172b", 
            x"13ec", x"0871", x"01e0", x"ffac", 
            x"f85d", x"f1e5", x"f08e", x"edd5", 
            x"e9f1", x"e920", x"eda2", x"f86c", 
            x"02d6", x"03d3", x"013c", x"04fc", 
            x"075b", x"fce9", x"eb08", x"deb1", 
            x"e008", x"ed0b", x"f619", x"ee4e", 
            x"e330", x"e8ea", x"f7fa", x"ff67", 
            x"ff1d", x"fe82", x"ff92", x"fcaf", 
            x"f65c", x"fa04", x"0715", x"09ad", 
            x"fe7b", x"f5e0", x"f26c", x"eee5", 
            x"f3f5", x"059f", x"1143", x"09bd", 
            x"fef2", x"01f4", x"0d54", x"1317", 
            x"0d44", x"02d6", x"fdd4", x"fed5", 
            x"fc44", x"f16f", x"ebf6", x"f492", 
            x"ffbf", x"055d", x"0407", x"fa6e", 
            x"ef3e", x"ed5a", x"f622", x"ff59", 
            x"ff19", x"f2a8", x"e551", x"e94f", 
            x"f98a", x"01f6", x"004e", x"fee5", 
            x"ff37", x"fbce", x"f7c5", x"fa84", 
            x"fecb", x"fdde", x"fdb5", x"01fa", 
            x"02e3", x"fc8a", x"f9e4", x"04ec", 
            x"1334", x"12bd", x"0559", x"f9c7", 
            x"f475", x"f412", x"fb6a", x"0a31", 
            x"1757", x"1a97", x"181e", x"17f2", 
            x"1760", x"136b", x"13c8", x"19eb", 
            x"19e0", x"10be", x"0c96", x"15a0", 
            x"20be", x"223a", x"1e29", x"1a31", 
            x"12cc", x"06b3", x"f93f", x"ec8f", 
            x"e473", x"e386", x"ea19", x"f5d5", 
            x"f8af", x"ebc8", x"e0ef", x"e49a", 
            x"ec3b", x"ef50", x"f154", x"f5bc", 
            x"f79e", x"f05c", x"ea6a", x"f09f", 
            x"f712", x"f2d9", x"eb34", x"e7dc", 
            x"e896", x"f007", x"0002", x"0ff4", 
            x"13bc", x"0c6d", x"0932", x"0ca4", 
            x"090e", x"fd83", x"f772", x"f92c", 
            x"fd34", x"03a7", x"0907", x"0c08", 
            x"14a9", x"2178", x"26a6", x"1d76", 
            x"0c29", x"02ee", x"02bf", x"fc43", 
            x"f261", x"f982", x"0f7d", x"1c69", 
            x"19ea", x"1153", x"065a", x"fbf3", 
            x"f607", x"f47c", x"f6ed", x"fedf", 
            x"0701", x"0bee", x"173c", x"2862", 
            x"2b86", x"1891", x"044f", x"0467", 
            x"0f52", x"0dbb", x"0684", x"0dde", 
            x"1b5b", x"19f3", x"0eb5", x"0ca7", 
            x"0e5c", x"044a", x"f5ac", x"f1bc", 
            x"f6a2", x"fb4c", x"fcd2", x"fcab", 
            x"f9d9", x"f0cd", x"e5c7", x"e856", 
            x"fc24", x"0a1d", x"019e", x"ef25", 
            x"e7d0", x"efa2", x"f8ff", x"f78f", 
            x"f1ce", x"f675", x"0347", x"0684", 
            x"fb55", x"f5c9", x"0652", x"1c7c", 
            x"1aff", x"0231", x"eebc", x"f59b", 
            x"0ca5", x"1667", x"0732", x"f1e8", 
            x"ee3f", x"fddd", x"08df", x"fe9e", 
            x"f271", x"fd97", x"116f", x"0c28", 
            x"f14d", x"e156", x"e19e", x"e2ce", 
            x"e2d3", x"e29a", x"e21f", x"e85b", 
            x"f8df", x"0b2a", x"1261", x"0da7", 
            x"05d7", x"fbf1", x"ee15", x"e4dc", 
            x"e718", x"eeb6", x"f254", x"f204", 
            x"f780", x"05a9", x"0e2b", x"04cc", 
            x"f48b", x"f173", x"fcf3", x"042e", 
            x"fb2d", x"edbc", x"e92e", x"e9d3", 
            x"ea6c", x"ef82", x"fa4c", x"006d", 
            x"f952", x"f092", x"f280", x"f82c", 
            x"fae5", x"ff88", x"08c2", x"0fdd", 
            x"0e27", x"0554", x"ff42", x"05d1", 
            x"1869", x"279b", x"24d6", x"1739", 
            x"12ef", x"1921", x"196d", x"10c5", 
            x"0d3a", x"13a4", x"148a", x"0680", 
            x"f95f", x"fcb1", x"0817", x"0d95", 
            x"08ab", x"f9da", x"ea70", x"e4da", 
            x"e379", x"dd84", x"d8e0", x"de54", 
            x"e896", x"ebe9", x"e93d", x"e508", 
            x"dded", x"db83", x"e744", x"f194", 
            x"e783", x"db9a", x"ea07", x"083c", 
            x"1823", x"157c", x"110b", x"16d5", 
            x"247d", x"2c5c", x"28d5", x"212c", 
            x"1ad5", x"18e2", x"1c73", x"2010", 
            x"1ec5", x"1bc3", x"1c97", x"1da6", 
            x"147d", x"ffcc", x"ea70", x"e1ae", 
            x"e634", x"e74f", x"dc02", x"d4d5", 
            x"df99", x"ef57", x"f817", x"fde0", 
            x"ff91", x"fb38", x"fb30", x"0334", 
            x"0914", x"069c", x"fc02", x"f32a", 
            x"fb7d", x"10dd", x"1e83", x"1b6f", 
            x"115f", x"0c4b", x"0e79", x"1113", 
            x"14a2", x"1e76", x"2339", x"16ed", 
            x"08af", x"0c21", x"14d7", x"0984", 
            x"f06a", x"e39b", x"e82b", x"f1b6", 
            x"f69e", x"f5d2", x"f4da", x"f8b2", 
            x"0564", x"1561", x"1803", x"0df1", 
            x"0909", x"0b7c", x"0ac3", x"0497", 
            x"fac3", x"f4fe", x"f8b7", x"fce6", 
            x"ff2b", x"0799", x"12a8", x"1599", 
            x"12e6", x"12d8", x"142e", x"118a", 
            x"0d3a", x"0d75", x"125d", x"1213", 
            x"0592", x"f955", x"ff6d", x"145f", 
            x"246d", x"26f7", x"20f1", x"1a0f", 
            x"15eb", x"0fab", x"0384", x"f8fd", 
            x"fabb", x"072d", x"0c27", x"0044", 
            x"f6e3", x"fea6", x"0929", x"0531", 
            x"fa70", x"f725", x"f60b", x"f6f5", 
            x"0583", x"14ae", x"0e24", x"fb96", 
            x"f31a", x"f84f", x"fe19", x"fd04", 
            x"ff66", x"08d0", x"0c44", x"049b", 
            x"fb78", x"fbdd", x"0316", x"0379", 
            x"01a6", x"0956", x"0f55", x"0e48", 
            x"11a7", x"14d7", x"0ea6", x"04bc", 
            x"fd7f", x"ff7c", x"07fe", x"035a", 
            x"f1a0", x"e693", x"e206", x"d974", 
            x"cddd", x"c793", x"cb5b", x"d36b", 
            x"da7f", x"e06f", x"e50a", x"e9bf"
        ),
        -- Block 9
        (
            x"ed96", x"eba0", x"e160", x"d4c4", 
            x"d3a2", x"e097", x"ece6", x"ef27", 
            x"ec1b", x"e9e1", x"ee9c", x"ff50", 
            x"1229", x"19a7", x"19a0", x"1ba5", 
            x"1ebe", x"1cbb", x"16ab", x"185e", 
            x"26e1", x"33c1", x"31ae", x"25c5", 
            x"1dd3", x"1f54", x"2146", x"19c9", 
            x"07e6", x"f5a3", x"eefc", x"f1ae", 
            x"f1b6", x"ebba", x"e80e", x"ea9c", 
            x"ec93", x"e7a7", x"db55", x"ce81", 
            x"ceaa", x"e035", x"f244", x"f34d", 
            x"e856", x"dfb2", x"e18c", x"ee1d", 
            x"fbc8", x"003d", x"ff03", x"03d3", 
            x"1016", x"1913", x"1be8", x"1fa2", 
            x"1fe9", x"181a", x"15db", x"1ec1", 
            x"1ec0", x"0d29", x"ff21", x"0424", 
            x"1178", x"14ad", x"0cc7", x"0adc", 
            x"12e7", x"1491", x"0a66", x"fcf5", 
            x"f2ec", x"f210", x"fd7f", x"0c6b", 
            x"0f8b", x"022b", x"eec8", x"e6dd", 
            x"f0ef", x"0143", x"08f8", x"0053", 
            x"ea6e", x"d9ba", x"e17d", x"fa57", 
            x"09f7", x"0a6b", x"0ae2", x"0959", 
            x"ff18", x"fac7", x"0564", x"0e89", 
            x"0863", x"fed6", x"ff4f", x"019f", 
            x"fdb4", x"fdf9", x"07f4", x"1035", 
            x"0d72", x"0437", x"fea7", x"0121", 
            x"03f6", x"fd23", x"f23f", x"f30f", 
            x"0216", x"0e6b", x"0e05", x"0a3c", 
            x"0816", x"04b2", x"0054", x"fb17", 
            x"f53b", x"f03f", x"eb95", x"e6cd", 
            x"e4f9", x"e814", x"f2e1", x"0069", 
            x"febb", x"eddb", x"e46c", x"ec5c", 
            x"fb01", x"04b0", x"0367", x"f8d5", 
            x"edeb", x"eccb", x"f7f7", x"0623", 
            x"0824", x"fcdc", x"f937", x"0625", 
            x"0c8d", x"fc5a", x"ec95", x"f6dd", 
            x"0dfe", x"15ae", x"0937", x"f93f", 
            x"f5dd", x"fd70", x"02d1", x"0272", 
            x"fd6c", x"f488", x"ee7a", x"f292", 
            x"ff90", x"0459", x"f3b5", x"dfaa", 
            x"dff8", x"ef95", x"faa3", x"f7fb", 
            x"f2de", x"f868", x"01c3", x"0180", 
            x"fa49", x"f976", x"0538", x"1405", 
            x"139e", x"0391", x"fc48", x"0dc8", 
            x"21aa", x"1931", x"016f", x"ffaa", 
            x"123f", x"17e3", x"0a9f", x"00d0", 
            x"010f", x"fbd5", x"f364", x"f9ef", 
            x"024f", x"f4dc", x"e48e", x"ed78", 
            x"ff70", x"ff39", x"f37a", x"f0e4", 
            x"f986", x"0398", x"0b6e", x"136a", 
            x"1c8e", x"2202", x"1d1d", x"0fa7", 
            x"0598", x"094a", x"1279", x"0f84", 
            x"0579", x"058d", x"0b90", x"057b", 
            x"f695", x"f21b", x"f674", x"f4da", 
            x"f0cb", x"f30e", x"f831", x"fcab", 
            x"0195", x"0659", x"064f", x"fd1c", 
            x"f0c9", x"ed25", x"f618", x"ff1a", 
            x"f8d7", x"e823", x"e542", x"fe39", 
            x"1c26", x"2097", x"1131", x"07b3", 
            x"076b", x"02b3", x"fa6e", x"f6a6", 
            x"f51c", x"f461", x"fb99", x"0e3f", 
            x"1fff", x"219c", x"12f5", x"0156", 
            x"fe31", x"0a39", x"0e9f", x"fbc7", 
            x"e471", x"e3be", x"f525", x"00d4", 
            x"ffff", x"ff5a", x"03ce", x"02ea", 
            x"f95d", x"f379", x"f8d9", x"01cf", 
            x"04b0", x"023f", x"fc3a", x"f27b", 
            x"f0f8", x"fd66", x"021d", x"f407", 
            x"e96d", x"ebbe", x"ea8a", x"e581", 
            x"e68b", x"e582", x"db60", x"d35c", 
            x"d4f5", x"dc96", x"e200", x"dbcc", 
            x"d097", x"d256", x"df5b", x"e7b3", 
            x"e858", x"eacc", x"f67d", x"056d", 
            x"088b", x"feaf", x"fbea", x"033a", 
            x"00f9", x"fb09", x"0856", x"1d5c", 
            x"2328", x"1f15", x"2101", x"2c35", 
            x"352b", x"2fe1", x"1a0a", x"0076", 
            x"fb0e", x"0e57", x"1edf", x"17ac", 
            x"04a1", x"fbf8", x"fd2f", x"f997", 
            x"f17c", x"ec35", x"e60e", x"df46", 
            x"e255", x"ed9b", x"f3f3", x"ee81", 
            x"e0ba", x"d969", x"e58b", x"f941", 
            x"011d", x"fe1d", x"fc27", x"02a2", 
            x"0802", x"fe45", x"f77e", x"0973", 
            x"1f43", x"225c", x"1da8", x"2064", 
            x"2bc9", x"36b9", x"3b54", x"3b6c", 
            x"2f6c", x"144f", x"0495", x"12ff", 
            x"29a3", x"3107", x"29a4", x"1b6f", 
            x"1631", x"2537", x"3794", x"3588", 
            x"2116", x"0ce9", x"01ed", x"fc7d", 
            x"f85c", x"f255", x"eb66", x"eb56", 
            x"f893", x"0b58", x"0f03", x"052e", 
            x"07f2", x"17cd", x"1ac7", x"0c0e", 
            x"fd77", x"f7d3", x"fa75", x"035c", 
            x"0880", x"00d2", x"f743", x"fd7c", 
            x"0f52", x"1da8", x"28f4", x"30b1", 
            x"2613", x"1105", x"0bdd", x"1787", 
            x"216a", x"1db4", x"13d2", x"1533", 
            x"1e7a", x"2153", x"1de4", x"127e", 
            x"fc9a", x"ed97", x"f54e", x"0461", 
            x"0326", x"f0bd", x"dfa9", x"db66", 
            x"de35", x"e561", x"efd7", x"f2a7", 
            x"ed87", x"ef34", x"f964", x"012a", 
            x"02c8", x"00fe", x"fa4f", x"f138", 
            x"ee74", x"f49b", x"fabd", x"f587", 
            x"ee00", x"f993", x"1711", x"2740", 
            x"1ab1", x"0c04", x"1001", x"1782", 
            x"1516", x"0d81", x"02a8", x"f8a4", 
            x"f5d4", x"f1d6", x"e695", x"dfee", 
            x"e2cd", x"e21e", x"d6c6", x"d050", 
            x"df5f", x"f619", x"fddb", x"f826", 
            x"ee7e", x"e4a9", x"e010", x"e5ca", 
            x"f27c", x"fabb", x"f962", x"fa0e", 
            x"0097", x"00b1", x"fb78", x"fb6e", 
            x"00c0", x"0181", x"f6a9", x"e8a3", 
            x"e9ec", x"fd35", x"0c3f", x"0c1b", 
            x"09bc", x"0bb5", x"0da8", x"0d39", 
            x"0722", x"fd64", x"fa71", x"ff3a", 
            x"ffa5", x"f48a", x"e588", x"e136", 
            x"eb8d", x"f158", x"e4b9", x"d4ea", 
            x"d347", x"d90c", x"de1d", x"ebb5", 
            x"fd47", x"0002", x"f2d1", x"e897", 
            x"ef0a", x"f66e", x"e999", x"d6b6", 
            x"d9ae", x"ee5f", x"fa2c", x"f4a6", 
            x"f157", x"fbda", x"040f", x"00eb", 
            x"006f", x"03ea", x"fcd2", x"ee43", 
            x"eaf4", x"faae", x"067c", x"f608", 
            x"deba", x"e040", x"f24d", x"fbc8", 
            x"f8b9", x"f4e6", x"ef6b", x"e47f", 
            x"e858", x"025c", x"11c5", x"0757", 
            x"f920", x"f5e3", x"f881", x"f672", 
            x"f44a", x"fe2f", x"0d68", x"12ac", 
            x"087c", x"f604", x"f274", x"08cb", 
            x"1cdc", x"1271", x"f852", x"f06c", 
            x"fc7e", x"0569", x"08f2", x"1133", 
            x"15aa", x"0c40", x"ffd0", x"fdcc", 
            x"fdf5", x"f4d3", x"ebdf", x"ee31", 
            x"f418", x"f535", x"f9f9", x"0466", 
            x"0641", x"00d4", x"ffda", x"fcb8", 
            x"eebc", x"e682", x"f478", x"064e", 
            x"08a4", x"0458", x"04d8", x"07c3", 
            x"0649", x"0119", x"ff02", x"fe51", 
            x"f8b4", x"f4cb", x"f9fc", x"037c", 
            x"0b4d", x"0f17", x"0ed7", x"0d2d", 
            x"0881", x"fe36", x"f552", x"fc26", 
            x"1892", x"32d5", x"2cde", x"1599", 
            x"1124", x"1d69", x"2377", x"2099", 
            x"1d9d", x"1fc8", x"2726", x"2a6b", 
            x"22df", x"1355", x"01e9", x"f958", 
            x"fde1", x"04e2", x"01a7", x"f2e6", 
            x"e769", x"ee27", x"ff71", x"0630", 
            x"ff78", x"fa70", x"01b2", x"10c7", 
            x"15e0", x"037e", x"ea60", x"ed29", 
            x"0ba8", x"1a5a", x"04ed", x"edfd", 
            x"f327", x"069d", x"1138", x"10d4", 
            x"1102", x"171d", x"1df8", x"20bc", 
            x"15e3", x"0287", x"0757", x"2240", 
            x"2ce7", x"2099", x"1864", x"1f4c", 
            x"1f31", x"0da9", x"03eb", x"0bbc", 
            x"0cab", x"042f", x"0386", x"0809", 
            x"0a58", x"0e4d", x"15c3", x"1b14", 
            x"1565", x"07c4", x"fc32", x"ef9d", 
            x"e690", x"f346", x"0bf6", x"0e7c", 
            x"f9c0", x"ed3d", x"f47b", x"ff9b", 
            x"0107", x"f93b", x"ef81", x"eaf6", 
            x"f00e", x"fa61", x"ff67", x"01e4", 
            x"0869", x"0854", x"ffb9", x"00d5", 
            x"083e", x"0116", x"f630", x"ffd6", 
            x"13ae", x"14ed", x"0247", x"fbc0", 
            x"0f82", x"1dc1", x"11fb", x"02d6", 
            x"0436", x"0e6d", x"11ed", x"0aa8", 
            x"fde9", x"f1cd", x"f258", x"0103", 
            x"0571", x"f368", x"e35a", x"e762", 
            x"ef56", x"eef5", x"ed5b", x"f071", 
            x"fa61", x"0ac4", x"1473", x"0852", 
            x"f2d7", x"f118", x"00f8", x"003b", 
            x"e4c9", x"cc74", x"d302", x"ef59", 
            x"0237", x"feaa", x"ef35", x"e79e", 
            x"f369", x"05e3", x"0cf3", x"0749", 
            x"fce4", x"f598", x"f6de", x"fc26", 
            x"fe00", x"ff90", x"0428", x"08e5", 
            x"0bfe", x"0bb3", x"02e6", x"f3cc", 
            x"ee50", x"fadd", x"06d7", x"ff1c", 
            x"f122", x"faaf", x"1a43", x"2231", 
            x"fac7", x"d3cf", x"dacb", x"f4ad", 
            x"f43c", x"e0f8", x"d9d2", x"dfb7", 
            x"e773", x"f24d", x"fe6f", x"ffae", 
            x"f4fd", x"ed80", x"ee5b", x"ef9b", 
            x"f0e6", x"f5d3", x"fe04", x"0ac0", 
            x"1339", x"07c6", x"f1a0", x"ebd4", 
            x"ff42", x"16e8", x"14a6", x"fa26", 
            x"ee23", x"fba0", x"030a", x"f9b6", 
            x"f5fa", x"fdb4", x"02b1", x"0517", 
            x"06b5", x"0005", x"f7ba", x"fad2", 
            x"0457", x"0ca2", x"14c1", x"1705", 
            x"07cc", x"efae", x"ec43", x"040a", 
            x"1745", x"10d2", x"03db", x"0a35", 
            x"1f06", x"2d9f", x"313b", x"3107", 
            x"2b70", x"1a87", x"0a68", x"0b6f", 
            x"1560", x"14a7", x"0910", x"046e", 
            x"0e5b", x"1b1c", x"1b0f", x"0b73", 
            x"f853", x"f0ff", x"f846", x"00ef", 
            x"f8a9", x"de07", x"cbfa", x"d562", 
            x"f08f", x"0b6b", x"186e", x"1304", 
            x"030d", x"f5db", x"f017", x"f4da", 
            x"0743", x"1687", x"0ff2", x"014d", 
            x"05c5", x"200d", x"33d6", x"29a9", 
            x"1107", x"0b8f", x"1e75", x"2940", 
            x"1a9e", x"0edf", x"1a7e", x"251f", 
            x"1a7b", x"0712", x"f632", x"edc5", 
            x"f44c", x"0167", x"0a3c", x"12db", 
            x"1d13", x"1a33", x"07d2", x"fe4f", 
            x"0c4e", x"1c35", x"1220", x"faef", 
            x"fc05", x"1650", x"2042", x"075a", 
            x"f396", x"0531", x"1c62", x"1381", 
            x"f87d", x"eec6", x"fe4a", x"0e24", 
            x"091a", x"f8fd", x"f389", x"fd23", 
            x"0c7f", x"1379", x"07af", x"f55d", 
            x"f585", x"08ec", x"141a", x"0a91", 
            x"fe64", x"0154", x"0a92", x"053a", 
            x"f201", x"e474", x"e283", x"e84b", 
            x"f86f", x"0ad4", x"0bc3", x"faa9", 
            x"ec81", x"eb21", x"ed15", x"e8b3", 
            x"e2cb", x"e21a", x"e36f", x"e62b", 
            x"ee42", x"f745", x"f447", x"e2e1", 
            x"dad0", x"eb17", x"f8d5", x"f10a", 
            x"e5a0", x"e3e6", x"e8dc", x"ef17", 
            x"ed4a", x"e248", x"d7cc", x"d34e", 
            x"d3dd", x"d8df", x"dfbd", x"e2ed", 
            x"e220", x"e134", x"e156", x"e2c2", 
            x"e99e", x"efdf", x"e9d3", x"e09e", 
            x"e05b", x"e1c8", x"e20c", x"e189", 
            x"d8aa", x"cc8e", x"cc95", x"d8c4", 
            x"e03f", x"dce2", x"dc03", x"e072", 
            x"e3fa", x"eea1", x"fd09", x"fc8b", 
            x"ee94", x"e868", x"f3cf", x"fd61", 
            x"eecf", x"d5ad", x"d104", x"e6a6", 
            x"fcc1", x"fc01", x"ea8c", x"e075", 
            x"e856", x"f073", x"e9c0", x"e045", 
            x"e396", x"e88b", x"de65", x"d89b", 
            x"f35a", x"1398", x"0b92", x"f06e", 
            x"f6a8", x"195e", x"2aec", x"203f", 
            x"1108", x"121b", x"2355", x"2b19", 
            x"19d4", x"071a", x"0c2e", x"1e21", 
            x"2417", x"1969", x"1217", x"17a9", 
            x"1650", x"097c", x"0966", x"14fb", 
            x"14b2", x"0ae9", x"0898", x"0fd5", 
            x"1825", x"1a58", x"1671", x"12ce", 
            x"10ef", x"0cc9", x"0312", x"f6ad", 
            x"ef6b", x"ef74", x"f57e", x"feee", 
            x"04df", x"0679", x"055b", x"0094", 
            x"fe88", x"03bb", x"0a4e", x"0b9f", 
            x"06c9", x"03d5", x"0b29", x"16e2", 
            x"1c0f", x"18c4", x"1349", x"1623", 
            x"1fd0", x"1fd3", x"114a", x"0230"
        ),
        -- Block 8
        (
            x"fe80", x"06a8", x"0df4", x"0943", 
            x"0647", x"0e15", x"0a18", x"f3d1", 
            x"ecdc", x"096c", x"2b6f", x"29f3", 
            x"0aa2", x"f84e", x"08eb", x"2517", 
            x"2cf2", x"231e", x"1fed", x"2629", 
            x"2981", x"25c7", x"1d30", x"1654", 
            x"1764", x"1c55", x"1abf", x"0ff2", 
            x"0325", x"0109", x"0cd9", x"1b4d", 
            x"25e2", x"2a90", x"227c", x"1119", 
            x"0886", x"0c90", x"0dd4", x"0765", 
            x"0217", x"00db", x"fd6a", x"fe66", 
            x"0e36", x"1c1f", x"0f45", x"ef76", 
            x"de44", x"e78d", x"f277", x"ecdd", 
            x"e76c", x"eeb6", x"f727", x"f7ba", 
            x"f7f3", x"ffd9", x"074d", x"0219", 
            x"f2ae", x"ea6d", x"ec12", x"eba7", 
            x"ea9a", x"efe0", x"f700", x"f686", 
            x"f4cd", x"fd44", x"09db", x"0c27", 
            x"081e", x"10f6", x"29e3", x"3d7f", 
            x"36e8", x"1db5", x"10fc", x"2034", 
            x"2ebf", x"2068", x"04eb", x"fb2b", 
            x"083e", x"1796", x"1895", x"1189", 
            x"0cde", x"02ee", x"efac", x"e50b", 
            x"ef80", x"fe8a", x"fe15", x"f663", 
            x"fc74", x"0cc4", x"1407", x"108e", 
            x"0f81", x"1179", x"0926", x"f98c", 
            x"f4d0", x"f95d", x"f8e8", x"f5d4", 
            x"f5fe", x"ed65", x"d95b", x"d36b", 
            x"e863", x"0018", x"ffb9", x"e7bc", 
            x"cfe2", x"cc58", x"dbd4", x"eddd", 
            x"ee6e", x"d932", x"c62c", x"cf93", 
            x"eab8", x"f714", x"ee69", x"e4d4", 
            x"e46d", x"e4ee", x"df19", x"d6a6", 
            x"d99c", x"f08a", x"0a0f", x"0947", 
            x"ee7c", x"ddc1", x"ee4a", x"0fe4", 
            x"1b7d", x"0018", x"dd9f", x"d723", 
            x"e61c", x"f6a4", x"00a5", x"03e9", 
            x"07c6", x"0dda", x"0dd7", x"105d", 
            x"2032", x"2b1c", x"2333", x"0de2", 
            x"f714", x"ed78", x"f16e", x"f56f", 
            x"f407", x"f297", x"f4bd", x"f539", 
            x"f1cb", x"f24b", x"f85f", x"fbe0", 
            x"f6b5", x"ebd9", x"e8c7", x"f4bf", 
            x"fe09", x"f2a9", x"e2dc", x"e8f1", 
            x"fc33", x"0323", x"f929", x"f104", 
            x"fce1", x"11d4", x"17bf", x"0a4d", 
            x"f62f", x"e6e2", x"e641", x"f550", 
            x"045f", x"08d5", x"06d3", x"fc8b", 
            x"e99e", x"e088", x"e77e", x"f516", 
            x"f945", x"e6d5", x"d38f", x"d857", 
            x"e878", x"f4cb", x"fe0f", x"fddd", 
            x"f21f", x"ea1f", x"f373", x"06f4", 
            x"0b42", x"fb95", x"faf5", x"139d", 
            x"20c9", x"1145", x"fdfe", x"fe05", 
            x"0d84", x"1d36", x"26b1", x"28ac", 
            x"20cf", x"14a7", x"0d98", x"106c", 
            x"1d9b", x"2a63", x"2426", x"11cc", 
            x"0c86", x"18a7", x"253f", x"1bec", 
            x"fc47", x"ea89", x"f90b", x"06df", 
            x"ff02", x"f102", x"ed67", x"f31c", 
            x"fa9f", x"0667", x"0efc", x"0463", 
            x"f07d", x"e996", x"ef86", x"f2ce", 
            x"eb52", x"ea04", x"ffb6", x"18ab", 
            x"1ab6", x"06dc", x"f1cb", x"f55e", 
            x"1557", x"2e74", x"2791", x"1018", 
            x"01d9", x"0b5d", x"1f2e", x"1c33", 
            x"0532", x"02af", x"1e38", x"338c", 
            x"2d2f", x"1ec0", x"19b5", x"1a59", 
            x"1bfc", x"1f5a", x"25a5", x"2522", 
            x"16cf", x"093a", x"0818", x"0b47", 
            x"09c2", x"04be", x"f86e", x"eb17", 
            x"f46b", x"0c20", x"11d2", x"005a", 
            x"ec7d", x"e88c", x"f264", x"fe69", 
            x"05a0", x"033c", x"f59e", x"e77f", 
            x"e4cd", x"ed1c", x"f742", x"f6f5", 
            x"f36a", x"fba6", x"0c1f", x"180a", 
            x"164e", x"0a08", x"fc84", x"f6d8", 
            x"fdbd", x"05ef", x"0085", x"ef73", 
            x"e709", x"fa22", x"1a3f", x"27e8", 
            x"21c4", x"17ac", x"0eb6", x"08e0", 
            x"09b1", x"0ff8", x"116a", x"01b7", 
            x"e970", x"e726", x"fa5f", x"fa4f", 
            x"e530", x"e5f7", x"fce3", x"fff4", 
            x"ea86", x"dd9c", x"df5d", x"dd14", 
            x"d8a0", x"e044", x"edae", x"f07d", 
            x"f071", x"ff13", x"1164", x"0f90", 
            x"02c9", x"067b", x"1215", x"0b7c", 
            x"fcb5", x"fcb5", x"032e", x"ff26", 
            x"fec2", x"0f2f", x"176d", x"0952", 
            x"0266", x"1405", x"2760", x"25ef", 
            x"124c", x"04e2", x"0ce0", x"1375", 
            x"047d", x"f15f", x"eeab", x"fb78", 
            x"0281", x"f30c", x"dde3", x"dbed", 
            x"e84a", x"ebb9", x"de43", x"d08d", 
            x"cf52", x"d451", x"d80a", x"d8d3", 
            x"d78c", x"dcc6", x"eafc", x"f4fb", 
            x"f107", x"ea87", x"f765", x"0e74", 
            x"0eef", x"fca9", x"f26c", x"f03c", 
            x"f3ed", x"0516", x"14d4", x"0cae", 
            x"f120", x"e287", x"f06f", x"042e", 
            x"0e18", x"121b", x"0bbe", x"fc87", 
            x"f3a8", x"f0c2", x"ebc2", x"ebb1", 
            x"f8af", x"0171", x"f2ca", x"e0ec", 
            x"e45e", x"ef0f", x"ee71", x"ec0e", 
            x"f263", x"f08e", x"dc7a", x"d7ef", 
            x"f9dd", x"1a98", x"11b7", x"f6e9", 
            x"eccf", x"f58f", x"0bd2", x"1c74", 
            x"1068", x"f715", x"f2b8", x"0b1e", 
            x"2895", x"2da9", x"1b47", x"090d", 
            x"0688", x"14dd", x"262a", x"26f3", 
            x"16be", x"04e1", x"fd6e", x"0484", 
            x"156f", x"27e3", x"2d85", x"1da9", 
            x"0b1f", x"0509", x"022b", x"0151", 
            x"082a", x"0b18", x"009a", x"f2b4", 
            x"f214", x"0059", x"0ce4", x"10c6", 
            x"0faf", x"0292", x"eba8", x"e3bf", 
            x"f26a", x"00e1", x"01c4", x"00f5", 
            x"096e", x"186c", x"22ee", x"2338", 
            x"1e4b", x"16bd", x"0da5", x"0968", 
            x"1073", x"1ccf", x"1998", x"ff8e", 
            x"efa6", x"0ad7", x"2e98", x"2662", 
            x"0712", x"008e", x"10c2", x"1c7e", 
            x"167e", x"ff7a", x"e9bb", x"e962", 
            x"f5d6", x"f9b6", x"f1f3", x"ee6e", 
            x"f722", x"fbd3", x"f8cc", x"03fc", 
            x"1772", x"135f", x"feb9", x"fc93", 
            x"0d2c", x"0fcb", x"fcc1", x"ede0", 
            x"ee34", x"f1c4", x"f5fb", x"fc47", 
            x"fd28", x"fb39", x"00f9", x"0af7", 
            x"06f4", x"f14b", x"e29c", x"e938", 
            x"f94e", x"034a", x"fb93", x"e960", 
            x"ec39", x"09fb", x"1b70", x"1256", 
            x"0953", x"0251", x"f3cc", x"f488", 
            x"112a", x"2769", x"1d03", x"0828", 
            x"0185", x"0457", x"0747", x"0c83", 
            x"1416", x"0c80", x"f797", x"f8a1", 
            x"126f", x"1aca", x"042d", x"f017", 
            x"f119", x"ee90", x"db8b", x"d6b7", 
            x"e619", x"eb72", x"e733", x"eecb", 
            x"fc6f", x"0370", x"0874", x"11f1", 
            x"1d35", x"1735", x"fa37", x"e596", 
            x"f143", x"0f9f", x"1efa", x"0f8e", 
            x"fb28", x"ffc4", x"1265", x"1c52", 
            x"1d5c", x"1bb2", x"14b5", x"068b", 
            x"f854", x"f578", x"04e4", x"172a", 
            x"13e2", x"fd73", x"f19d", x"fec2", 
            x"0627", x"f549", x"e856", x"e7ba", 
            x"e066", x"d962", x"e00b", x"e754", 
            x"e15e", x"daca", x"e759", x"f94b", 
            x"f856", x"f220", x"f5b7", x"f33e", 
            x"e429", x"dcb4", x"eadb", x"0092", 
            x"0a02", x"043e", x"fe19", x"0119", 
            x"06fd", x"0c58", x"0ad1", x"fba9", 
            x"eba2", x"ecfb", x"f83b", x"fc69", 
            x"f9a9", x"f6ef", x"f6f3", x"0267", 
            x"19e3", x"1f69", x"0a32", x"fbb6", 
            x"02da", x"0c85", x"0c41", x"0c67", 
            x"0dd3", x"019c", x"f363", x"fca8", 
            x"0ba7", x"045a", x"f9ac", x"0048", 
            x"0cdd", x"115d", x"0c74", x"0447", 
            x"0013", x"00f2", x"029e", x"011c", 
            x"fba9", x"f747", x"fad5", x"02cf", 
            x"00c0", x"f6c8", x"f696", x"fc36", 
            x"f2a9", x"e06c", x"e08b", x"f0ed", 
            x"f5f8", x"ea05", x"e182", x"ec07", 
            x"03e4", x"1381", x"09db", x"f4dc", 
            x"f14e", x"ff8a", x"0b1c", x"0951", 
            x"ff70", x"facd", x"0684", x"1450", 
            x"0f4c", x"02f7", x"0759", x"1b4f", 
            x"25ed", x"1292", x"f093", x"eb95", 
            x"0b75", x"21da", x"0a54", x"ebb7", 
            x"f1d0", x"043e", x"0427", x"f779", 
            x"edd1", x"eabe", x"ee08", x"f810", 
            x"0176", x"f6c1", x"e18e", x"e599", 
            x"fcbb", x"01b0", x"f1aa", x"e7dc", 
            x"f22b", x"006b", x"0398", x"016a", 
            x"fe37", x"fd22", x"0884", x"1773", 
            x"1aab", x"1b09", x"1db5", x"1a7c", 
            x"14d5", x"121e", x"0998", x"015f", 
            x"0aef", x"2210", x"2b86", x"1719", 
            x"f65b", x"e869", x"f273", x"f868", 
            x"ea07", x"e176", x"f3aa", x"07bd", 
            x"040e", x"f836", x"fbfc", x"0db0", 
            x"1c64", x"1963", x"01fe", x"ea77", 
            x"ed5a", x"ffa1", x"02da", x"ff50", 
            x"0b32", x"121d", x"06e7", x"02a8", 
            x"0ba1", x"1210", x"15b1", x"19d2", 
            x"19cf", x"17f9", x"13b4", x"0b14", 
            x"01e4", x"f37c", x"e3bb", x"e4b1", 
            x"efbf", x"eeea", x"e3c3", x"e572", 
            x"fe2f", x"1392", x"11ce", x"0656", 
            x"fe48", x"fa96", x"f8b9", x"f155", 
            x"e441", x"e174", x"eb77", x"f5c7", 
            x"00c9", x"09b8", x"05de", x"0019", 
            x"faf9", x"ed65", x"ebdb", x"05dd", 
            x"20f1", x"24c5", x"209b", x"22c1", 
            x"1fe4", x"1900", x"17ba", x"14d2", 
            x"0aec", x"ff8e", x"fbe0", x"0106", 
            x"027c", x"fbfa", x"f79e", x"f512", 
            x"f3d7", x"fdf1", x"02a9", x"ecc8", 
            x"dd3e", x"f4e0", x"11e7", x"0cde", 
            x"f3ae", x"eac6", x"f4ac", x"ee0d", 
            x"d2de", x"ccc9", x"e402", x"f28e", 
            x"f387", x"0030", x"0b3f", x"fca7", 
            x"ee0d", x"f3a0", x"f5e0", x"ef82", 
            x"ed3a", x"f20c", x"fa3c", x"f767", 
            x"e7f6", x"e661", x"01ed", x"1d7b", 
            x"177a", x"fcec", x"f45b", x"01ac", 
            x"0ae9", x"0107", x"ee15", x"e4e2", 
            x"e41d", x"e442", x"ec35", x"f80b", 
            x"f51a", x"efe9", x"00c5", x"18c9", 
            x"14b2", x"f8a8", x"f45e", x"1496", 
            x"2ddf", x"22f3", x"02fa", x"f019", 
            x"febe", x"19a5", x"1d6e", x"0836", 
            x"f73d", x"f7ed", x"f7ea", x"ef3c", 
            x"ef36", x"0354", x"19e8", x"1c61", 
            x"0efc", x"076b", x"140e", x"2c4b", 
            x"3305", x"1baf", x"0633", x"0df3", 
            x"16a3", x"0218", x"f0ca", x"00e4", 
            x"0ed9", x"0227", x"fa2a", x"0226", 
            x"043b", x"0330", x"0a05", x"120d", 
            x"137a", x"1094", x"14d9", x"1c25", 
            x"1210", x"f9d0", x"ef67", x"fcb5", 
            x"0fe8", x"12d6", x"03d3", x"f40a", 
            x"f3ed", x"084e", x"1be7", x"141f", 
            x"01f9", x"000e", x"fd69", x"e8d0", 
            x"d6c7", x"e2b8", x"06f7", x"23b8", 
            x"1fd6", x"02e0", x"f535", x"0f86", 
            x"30d0", x"2c1f", x"0967", x"ed38", 
            x"e88b", x"f6c9", x"09d5", x"12d3", 
            x"0ad0", x"fbfb", x"f739", x"fc52", 
            x"0265", x"0b48", x"0fe6", x"04b1", 
            x"f66a", x"f74f", x"07cd", x"1067", 
            x"fadd", x"e0cb", x"ea09", x"02ef", 
            x"fea6", x"e611", x"e5d6", x"ff75", 
            x"0e69", x"0952", x"02a0", x"0058", 
            x"fe44", x"052e", x"15a6", x"18d3", 
            x"0825", x"fca9", x"060f", x"1769", 
            x"13c6", x"f807", x"e553", x"f6f9", 
            x"19a9", x"236f", x"0f26", x"f769", 
            x"f1e9", x"fa1b", x"fdca", x"f64a", 
            x"e9e1", x"dc33", x"d4a1", x"daaf", 
            x"de02", x"ce46", x"b6b0", x"af1a", 
            x"c141", x"d608", x"d61e", x"cddd", 
            x"cea2", x"da99", x"ecb4", x"fb35", 
            x"f87b", x"e421", x"d8f6", x"ec90", 
            x"08d2", x"0887", x"f8a3", x"0719", 
            x"2b9f", x"33e0", x"2351", x"20d8", 
            x"2582", x"1c4e", x"14a6", x"1cc4", 
            x"1d30", x"0618", x"f081", x"ee61", 
            x"ef54", x"e3b6", x"d54b", x"cf42", 
            x"cd47", x"cb70", x"d4dc", x"e5a4", 
            x"e4d1", x"d234", x"c965", x"d5cf", 
            x"e49a", x"e779", x"e77e", x"e71b", 
            x"de37", x"d943", x"e789", x"f6a2", 
            x"f72f", x"fd51", x"1614", x"263c"
        ),
        -- Block 7
        (
            x"17a8", x"0a34", x"1cf4", x"328c", 
            x"2ced", x"1d9f", x"141a", x"0848", 
            x"04ca", x"1f7c", x"3aa4", x"2751", 
            x"fe75", x"f406", x"fe63", x"f631", 
            x"de31", x"d75f", x"e5d4", x"f2af", 
            x"fab6", x"0948", x"0db0", x"029e", 
            x"06f1", x"18e2", x"144d", x"fb6f", 
            x"efb2", x"f8df", x"03c8", x"0301", 
            x"0423", x"109a", x"156f", x"079e", 
            x"feff", x"0e12", x"2703", x"2c1e", 
            x"1b7b", x"112e", x"141e", x"12de", 
            x"07e2", x"0192", x"05a0", x"04ca", 
            x"fae1", x"f6cb", x"fa48", x"fe61", 
            x"fee2", x"ffd7", x"0549", x"0437", 
            x"f8be", x"f599", x"ffd7", x"0028", 
            x"efde", x"e874", x"fa2b", x"0e58", 
            x"0d8e", x"0089", x"fb8a", x"0434", 
            x"123f", x"1ce4", x"1d92", x"0ffb", 
            x"011e", x"0035", x"0654", x"0bc8", 
            x"1059", x"0f2c", x"0d8f", x"0bc2", 
            x"05c3", x"08ef", x"1133", x"146c", 
            x"1ccb", x"24d0", x"1113", x"edc2", 
            x"e9a8", x"05cd", x"138f", x"ffff", 
            x"ec3f", x"edcf", x"fda5", x"1a34", 
            x"33b7", x"2c73", x"0fdd", x"fe50", 
            x"fa32", x"f686", x"efa8", x"f259", 
            x"029b", x"08ff", x"03fb", x"04d6", 
            x"fe08", x"efc0", x"f9a5", x"14a0", 
            x"154c", x"f910", x"e656", x"ede8", 
            x"f6d7", x"f569", x"f7f3", x"f970", 
            x"f064", x"efd8", x"05fd", x"1c5d", 
            x"1bd3", x"1104", x"0d65", x"1086", 
            x"1865", x"2312", x"271f", x"1950", 
            x"00a5", x"f5ae", x"fd44", x"02df", 
            x"0039", x"ffb5", x"0068", x"fbf3", 
            x"f7cf", x"f915", x"f674", x"eeae", 
            x"e9e4", x"e917", x"ed8b", x"f6d2", 
            x"f9cf", x"f063", x"ea97", x"f3cd", 
            x"fd8f", x"fb4a", x"f501", x"ee52", 
            x"def3", x"d10c", x"dbab", x"f7be", 
            x"06a9", x"027a", x"fce9", x"fdb3", 
            x"01dd", x"062f", x"09d6", x"04ca", 
            x"faa3", x"01f9", x"124c", x"0ae4", 
            x"f432", x"ede7", x"f6be", x"fd1a", 
            x"01ea", x"0f47", x"167d", x"0675", 
            x"f230", x"f61a", x"053c", x"057d", 
            x"fb80", x"f1b2", x"f2e4", x"09f5", 
            x"229b", x"27e2", x"1d6f", x"0a69", 
            x"0718", x"1291", x"0c03", x"fdda", 
            x"ff03", x"003f", x"fd31", x"084e", 
            x"1428", x"1637", x"185b", x"1adf", 
            x"17ac", x"10ee", x"1402", x"171f", 
            x"10ad", x"0f5b", x"0df7", x"0340", 
            x"01a1", x"0747", x"08b6", x"0c56", 
            x"0b54", x"fea1", x"f079", x"ee0b", 
            x"fb66", x"0cbd", x"1455", x"0ffc", 
            x"0641", x"0506", x"0ddd", x"0c67", 
            x"0314", x"0761", x"104f", x"100e", 
            x"1275", x"18ac", x"1263", x"032e", 
            x"fd2e", x"0487", x"04d6", x"fa41", 
            x"fcd3", x"1095", x"20ab", x"1a22", 
            x"0807", x"0b68", x"1f25", x"1c54", 
            x"07ea", x"0308", x"0f98", x"1968", 
            x"1143", x"ffd0", x"ffc8", x"0985", 
            x"fc60", x"e372", x"e8a3", x"0f32", 
            x"3098", x"2ac1", x"08ee", x"f97d", 
            x"06b6", x"0e92", x"fd9e", x"eb2f", 
            x"f1e0", x"026e", x"015d", x"f4ba", 
            x"fafc", x"14fa", x"1e73", x"117b", 
            x"074d", x"fd65", x"f023", x"f3aa", 
            x"075d", x"0d84", x"ff1f", x"f44f", 
            x"f010", x"ed2e", x"f67a", x"fbaf", 
            x"e3bd", x"c76b", x"cafc", x"e1a8", 
            x"ec7c", x"e78a", x"e36a", x"e866", 
            x"eb2c", x"ea6a", x"f8a5", x"0df7", 
            x"0716", x"f00b", x"fb71", x"1e9b", 
            x"2a51", x"235a", x"1e9f", x"1193", 
            x"fe16", x"f810", x"ffa1", x"0472", 
            x"fd00", x"f38f", x"f41d", x"f8c3", 
            x"0217", x"0d1c", x"041c", x"e914", 
            x"dc59", x"e42d", x"e831", x"e111", 
            x"de6c", x"e6ec", x"e86c", x"daad", 
            x"d9c7", x"f47f", x"fbec", x"d876", 
            x"c72d", x"e8ad", x"01f5", x"e356", 
            x"b42e", x"af3e", x"d44f", x"f470", 
            x"ec08", x"d1be", x"cd93", x"e874", 
            x"0d7b", x"1d9f", x"12b0", x"0385", 
            x"fa04", x"f374", x"f7aa", x"013c", 
            x"1055", x"2a29", x"311a", x"1c2d", 
            x"0933", x"f828", x"f297", x"0c08", 
            x"1a77", x"f983", x"d267", x"d9eb", 
            x"fe09", x"0d9d", x"049e", x"f5ff", 
            x"e7c6", x"dfb9", x"de94", x"e128", 
            x"e9ab", x"ef57", x"e597", x"d7c0", 
            x"d1b0", x"d25a", x"e0ec", x"f34b", 
            x"f8f6", x"fdc0", x"0bb7", x"1253", 
            x"0199", x"ea4d", x"e67a", x"f4dd", 
            x"ff39", x"f846", x"edca", x"f112", 
            x"00e7", x"0f27", x"0c90", x"fa19", 
            x"ecf4", x"f6f0", x"06de", x"fec1", 
            x"e4d2", x"df66", x"0415", x"2e75", 
            x"2723", x"faaa", x"ea98", x"00b0", 
            x"0f7e", x"05dd", x"f9dc", x"f6c5", 
            x"ef0a", x"e8c9", x"f702", x"0bd4", 
            x"0aee", x"fa64", x"fafd", x"0c99", 
            x"0cf0", x"f8f2", x"ec24", x"f695", 
            x"10d4", x"2079", x"14e0", x"0038", 
            x"fe81", x"160f", x"3087", x"2fb1", 
            x"13d9", x"0300", x"1450", x"3078", 
            x"3276", x"0f8d", x"e99f", x"ed6c", 
            x"1159", x"1d2a", x"fba9", x"d7c4", 
            x"df49", x"025b", x"0b59", x"f70c", 
            x"ee7e", x"f049", x"e279", x"d788", 
            x"ebc6", x"ff94", x"eb47", x"d73b", 
            x"ee37", x"0938", x"ffbf", x"ed8e", 
            x"fb43", x"20b2", x"2af6", x"0cd7", 
            x"f72a", x"0095", x"0bde", x"0b5e", 
            x"0f4d", x"1826", x"1f8b", x"292c", 
            x"34dc", x"4048", x"3c22", x"2547", 
            x"18c0", x"1a61", x"1985", x"1b90", 
            x"1e6b", x"0e6f", x"fc0c", x"0565", 
            x"1d47", x"2329", x"0cb6", x"eabe", 
            x"d8cf", x"e0e6", x"f357", x"fd4a", 
            x"f726", x"e97f", x"e705", x"f513", 
            x"fef9", x"f4d6", x"e9c7", x"f8d9", 
            x"18c3", x"2b61", x"2f79", x"2d35", 
            x"263d", x"25e3", x"2b8d", x"2846", 
            x"1b3a", x"12d6", x"124a", x"1196", 
            x"11a5", x"0f8c", x"0a79", x"12a0", 
            x"22c5", x"24a3", x"1b34", x"10d0", 
            x"0806", x"0319", x"fc75", x"eef0", 
            x"e2d0", x"ddd2", x"e1af", x"ee6c", 
            x"f70e", x"f525", x"f264", x"f1e3", 
            x"f13f", x"f387", x"fb8e", x"042a", 
            x"fea4", x"edf6", x"eebe", x"08d2", 
            x"15c1", x"fe17", x"e653", x"f412", 
            x"104c", x"13f1", x"fe89", x"edab", 
            x"f4f5", x"0b6d", x"1aed", x"0a3b", 
            x"ec71", x"ea47", x"f787", x"fb05", 
            x"fd71", x"01db", x"000f", x"f44c", 
            x"e27c", x"dcd1", x"ed50", x"fa4a", 
            x"f09d", x"e5c9", x"ed82", x"0094", 
            x"0844", x"0276", x"f96c", x"efb9", 
            x"fa2c", x"1bf5", x"270a", x"0796", 
            x"df32", x"d38b", x"f340", x"1d68", 
            x"1585", x"e1e0", x"cf6a", x"f29d", 
            x"07d0", x"efe3", x"e23d", x"f5b6", 
            x"f648", x"dbfc", x"de74", x"006f", 
            x"1205", x"0187", x"e571", x"e0fa", 
            x"f1f3", x"fcf3", x"0394", x"0795", 
            x"fe11", x"f149", x"f8a7", x"100a", 
            x"19dc", x"0ba7", x"fd67", x"fc1f", 
            x"fff7", x"ffd8", x"f873", x"f2d4", 
            x"f8bc", x"02e4", x"feee", x"f448", 
            x"ffa7", x"15e7", x"0db9", x"f871", 
            x"fce2", x"0839", x"0607", x"05a3", 
            x"0a5b", x"05f7", x"fb56", x"f623", 
            x"f841", x"fb9e", x"f5d5", x"eb72", 
            x"e819", x"ebba", x"f131", x"f9b2", 
            x"06d3", x"19cc", x"2848", x"1cce", 
            x"0266", x"fff9", x"1a7c", x"21b0", 
            x"061b", x"f432", x"fd5f", x"046e", 
            x"f756", x"eb10", x"f67b", x"0fc2", 
            x"1b71", x"165a", x"0fc8", x"056e", 
            x"fd78", x"08f5", x"143a", x"07c5", 
            x"f560", x"f271", x"f82d", x"017a", 
            x"1022", x"137f", x"03a0", x"001b", 
            x"1ae1", x"3144", x"2930", x"14d7", 
            x"0c81", x"16a0", x"25fc", x"1f06", 
            x"fe2f", x"e722", x"eafb", x"fb05", 
            x"0b7a", x"1199", x"0bdd", x"0822", 
            x"0ea4", x"19ae", x"1fb9", x"1100", 
            x"ee48", x"da4e", x"e78d", x"f600", 
            x"ef50", x"e60f", x"e294", x"e431", 
            x"f25e", x"0847", x"1731", x"0ee0", 
            x"ee7a", x"d8da", x"eb10", x"0aa5", 
            x"0b1f", x"f612", x"f96b", x"17fa", 
            x"2478", x"0e39", x"fb0d", x"01b6", 
            x"0b58", x"fb36", x"e494", x"fc01", 
            x"3286", x"41a0", x"1733", x"e9b5", 
            x"e97e", x"0e77", x"2e88", x"2a05", 
            x"0174", x"e122", x"eccd", x"01a9", 
            x"fad0", x"e7b3", x"df03", x"e1c6", 
            x"eb08", x"f44d", x"f84a", x"f21d", 
            x"e547", x"e343", x"fa99", x"12b1", 
            x"0655", x"ec7c", x"eed2", x"09ea", 
            x"226d", x"1fe3", x"0758", x"fed2", 
            x"0bdd", x"0b64", x"fc29", x"0117", 
            x"1015", x"0476", x"efe5", x"f2f3", 
            x"fcf7", x"f9e6", x"f88e", x"f96c", 
            x"e843", x"daff", x"eca5", x"fd5b", 
            x"f1d9", x"e1cb", x"e044", x"e7ef", 
            x"ea32", x"e154", x"e929", x"021f", 
            x"0b7e", x"098e", x"0786", x"f685", 
            x"ed98", x"0def", x"286f", x"07cc", 
            x"d853", x"d9c0", x"f90c", x"04e3", 
            x"fce2", x"f5f7", x"ef7a", x"eb30", 
            x"f1cc", x"0949", x"2542", x"21e3", 
            x"0491", x"f628", x"fb2f", x"fbd0", 
            x"eda7", x"dae4", x"dbe0", x"ef7f", 
            x"fcea", x"fe10", x"fffb", x"0eb4", 
            x"177e", x"08f1", x"fd63", x"0464", 
            x"033f", x"fa7b", x"fc8e", x"fbbb", 
            x"f1fd", x"f6df", x"14d8", x"21e2", 
            x"0a0b", x"fa29", x"05be", x"115c", 
            x"1528", x"13f8", x"fd9c", x"e99b", 
            x"fc22", x"1719", x"0d86", x"f013", 
            x"f175", x"1175", x"1fe4", x"0854", 
            x"e88d", x"e8b4", x"0871", x"1c7b", 
            x"0cc4", x"f81e", x"f7ed", x"f92e", 
            x"f8ad", x"07cd", x"1947", x"18ab", 
            x"1000", x"0afd", x"07f3", x"0ccf", 
            x"1bc1", x"2519", x"1b0f", x"0420", 
            x"f1bf", x"f457", x"0544", x"10c2", 
            x"0f7e", x"0a6e", x"0660", x"0230", 
            x"0232", x"0565", x"03a0", x"f964", 
            x"f181", x"f5d0", x"0092", x"fdc5", 
            x"edf6", x"ed11", x"fb89", x"f800", 
            x"df8f", x"d321", x"e200", x"f056", 
            x"e94d", x"e2e3", x"f7c2", x"1aae", 
            x"2345", x"05d8", x"df80", x"cf47", 
            x"e331", x"030b", x"0013", x"e350", 
            x"dfc5", x"f52e", x"083a", x"1f8c", 
            x"2c81", x"0ab4", x"d7b9", x"d7b9", 
            x"04b1", x"181b", x"ff71", x"eefa", 
            x"003e", x"13d4", x"1403", x"1286", 
            x"1d69", x"1cf2", x"03d9", x"f26a", 
            x"fff0", x"198e", x"1da2", x"08cf", 
            x"03dd", x"1bea", x"2b2e", x"1481", 
            x"f14b", x"f13e", x"0fa5", x"17fc", 
            x"01c3", x"f7a8", x"fdbb", x"fd35", 
            x"f89f", x"0504", x"16d4", x"1432", 
            x"03e4", x"fc32", x"ffec", x"0fb4", 
            x"1f07", x"1402", x"feba", x"0292", 
            x"1aa1", x"1cd4", x"f650", x"d635", 
            x"e84e", x"0d40", x"106f", x"f683", 
            x"eb67", x"f61c", x"fd12", x"fa82", 
            x"f158", x"e041", x"d6af", x"e74d", 
            x"0635", x"136a", x"05ff", x"f928", 
            x"fd13", x"074e", x"1921", x"311d", 
            x"35d1", x"1c4b", x"0002", x"07af", 
            x"23a6", x"19f3", x"f246", x"e6e6", 
            x"fddc", x"158f", x"1366", x"0374", 
            x"051e", x"162a", x"1de3", x"0f8d", 
            x"fa62", x"eb4e", x"e4ee", x"ed38", 
            x"0277", x"057a", x"e75f", x"d4cb", 
            x"f38c", x"16ff", x"00af", x"d138", 
            x"d26d", x"febf", x"0aca", x"e5f6", 
            x"d54c", x"ed31", x"0263", x"0b24", 
            x"1109", x"0ef5", x"0af4", x"1078", 
            x"1a2a", x"1abb", x"0b7d", x"012f", 
            x"095a", x"0b2d", x"ff18", x"fc7a", 
            x"1356", x"28cb", x"15c5", x"eebc", 
            x"e46b", x"f130", x"f7f3", x"f86e", 
            x"f061", x"e4c2", x"e1fc", x"e481", 
            x"ea6b", x"f17b", x"f143", x"edfb"
        ),
        -- Block 6
        (
            x"f36c", x"04eb", x"1bd3", x"1dd7", 
            x"ff66", x"e87f", x"f482", x"0547", 
            x"06ff", x"01cd", x"fff5", x"0d53", 
            x"1b79", x"110c", x"ff70", x"0ff5", 
            x"28a0", x"1084", x"e75d", x"ee7d", 
            x"0cb8", x"0926", x"edf7", x"ecd2", 
            x"12e2", x"29bb", x"0e39", x"eec9", 
            x"ee33", x"f13f", x"e675", x"e49d", 
            x"eeb2", x"e875", x"d0c5", x"c46e", 
            x"ce19", x"e410", x"f742", x"f307", 
            x"e69f", x"f194", x"014c", x"fe95", 
            x"f737", x"f5ac", x"f399", x"ed00", 
            x"ed33", x"f68f", x"fdb1", x"06af", 
            x"1b23", x"2470", x"1981", x"19e2", 
            x"2cda", x"2cb7", x"03ac", x"df8b", 
            x"edb0", x"0d40", x"107b", x"05ac", 
            x"0022", x"f93a", x"ee9b", x"e7d5", 
            x"e9a7", x"e198", x"cdfd", x"ccd5", 
            x"d96b", x"d62f", x"c84b", x"c638", 
            x"d2da", x"e3b4", x"ec82", x"ed10", 
            x"e915", x"e7a9", x"ee7b", x"f227", 
            x"ec00", x"f122", x"0982", x"1a33", 
            x"24ce", x"318c", x"25eb", x"03c6", 
            x"f6d8", x"0a52", x"17fe", x"0f44", 
            x"0771", x"0a4e", x"08b9", x"0324", 
            x"096f", x"1222", x"0d99", x"053e", 
            x"0536", x"04a2", x"f788", x"ec87", 
            x"f35f", x"01d8", x"0a08", x"038f", 
            x"f938", x"00d8", x"0bb2", x"0095", 
            x"eba3", x"e474", x"f476", x"0be6", 
            x"06f1", x"ee33", x"f73b", x"1ded", 
            x"2758", x"1016", x"08be", x"10d2", 
            x"0481", x"f778", x"ff4a", x"ff9f", 
            x"f1c7", x"f65c", x"1545", x"3283", 
            x"2d2b", x"0783", x"f316", x"0901", 
            x"1f2b", x"13ad", x"ff0b", x"09a6", 
            x"2bf1", x"325a", x"1e06", x"1a3f", 
            x"1fda", x"1162", x"fad6", x"f6a3", 
            x"0056", x"0a30", x"0d93", x"1061", 
            x"18b3", x"14d4", x"fe7e", x"ee59", 
            x"f9a2", x"0cdf", x"0d0c", x"ff54", 
            x"0218", x"1435", x"0af2", x"f1d9", 
            x"fcca", x"14ae", x"13eb", x"0772", 
            x"fefe", x"0196", x"047a", x"feb9", 
            x"0315", x"0e7b", x"0605", x"fd4c", 
            x"0fb7", x"23c2", x"249a", x"15bd", 
            x"0c6f", x"153e", x"18eb", x"103c", 
            x"0c4e", x"103c", x"1363", x"1496", 
            x"151b", x"1aa8", x"1ea7", x"176a", 
            x"0791", x"f224", x"e940", x"facd", 
            x"08de", x"f9f6", x"ea01", x"f4bb", 
            x"08c7", x"08e4", x"f53d", x"f46f", 
            x"1117", x"1dd7", x"107f", x"075a", 
            x"05f3", x"0343", x"0182", x"0751", 
            x"1a19", x"23e0", x"18a6", x"1253", 
            x"09bb", x"f3cf", x"ebd2", x"f4e5", 
            x"f7ef", x"f570", x"f31d", x"e87e", 
            x"df3e", x"e334", x"f47d", x"0c0b", 
            x"0bc6", x"ec3f", x"df46", x"fbcc", 
            x"1f41", x"2c7b", x"26d8", x"1608", 
            x"07dc", x"11c4", x"231b", x"14df", 
            x"f12f", x"e424", x"f4d9", x"0496", 
            x"0071", x"fb8e", x"0c62", x"222e", 
            x"2566", x"13f3", x"fd4a", x"f1dc", 
            x"ef1a", x"eda9", x"e019", x"c1a6", 
            x"bd72", x"e409", x"00de", x"fa21", 
            x"ef7c", x"f41d", x"f5d9", x"ea82", 
            x"d657", x"d0d6", x"e8c4", x"0642", 
            x"0a6a", x"f96e", x"e898", x"e6d1", 
            x"f0ed", x"0016", x"15b6", x"1ba3", 
            x"0bef", x"0b7b", x"175d", x"1246", 
            x"01ca", x"f93f", x"ff81", x"08ba", 
            x"f7f9", x"da89", x"de0c", x"f66c", 
            x"0773", x"11c9", x"0e19", x"fcd8", 
            x"f70c", x"0046", x"0155", x"f5ef", 
            x"ee13", x"e996", x"e5d0", x"eab8", 
            x"ec27", x"dfa8", x"e1b8", x"f727", 
            x"028a", x"fda4", x"f160", x"e91f", 
            x"f444", x"0396", x"f8ed", x"e6b4", 
            x"e17e", x"e67d", x"fe57", x"104d", 
            x"01d5", x"e85d", x"d9be", x"e448", 
            x"fd37", x"fa99", x"e602", x"e7c1", 
            x"fc0b", x"00c1", x"e8f7", x"d942", 
            x"e219", x"e854", x"e606", x"e15f", 
            x"d9da", x"dfe8", x"ee3c", x"ed6b", 
            x"ec70", x"f6ff", x"f6f4", x"f153", 
            x"f86b", x"ff69", x"0a68", x"23dd", 
            x"31cd", x"1fb5", x"04d6", x"fccf", 
            x"0399", x"0c7e", x"120d", x"14c5", 
            x"1814", x"1667", x"07b2", x"fada", 
            x"04ee", x"15da", x"0b10", x"f2d6", 
            x"f2ea", x"01ad", x"05a6", x"0094", 
            x"f8c5", x"f2b8", x"f559", x"fe6e", 
            x"ff2c", x"f62f", x"f43f", x"f3f3", 
            x"ecfd", x"dd87", x"d0d8", x"e9f7", 
            x"2358", x"3635", x"14f6", x"06e3", 
            x"1cac", x"2c6b", x"281e", x"198e", 
            x"06d7", x"f3b7", x"ecdf", x"f79c", 
            x"05e7", x"068f", x"f4b8", x"e6c1", 
            x"f62a", x"1261", x"1b9e", x"1458", 
            x"0ca3", x"07a9", x"02ff", x"004e", 
            x"0642", x"15e3", x"15f6", x"ff8f", 
            x"f401", x"0329", x"1b8c", x"276e", 
            x"1bc4", x"0a2c", x"12bb", x"2bca", 
            x"34b8", x"288d", x"1a99", x"1cee", 
            x"234b", x"17b4", x"0e15", x"15bd", 
            x"1bda", x"153b", x"055a", x"f3bd", 
            x"eecf", x"f7d2", x"0728", x"0c13", 
            x"fc06", x"e8ce", x"e3a9", x"f29e", 
            x"0904", x"033c", x"dfde", x"cf75", 
            x"d63a", x"d75d", x"d0d5", x"c3c5", 
            x"bd0c", x"c82f", x"e0cc", x"f9cf", 
            x"f604", x"e19f", x"e0f8", x"e340", 
            x"dcb9", x"dcc6", x"e012", x"df9b", 
            x"eb39", x"0f15", x"3324", x"372d", 
            x"1c49", x"0578", x"0281", x"fc68", 
            x"e6fb", x"d81b", x"e46c", x"ffb1", 
            x"0952", x"fbad", x"f593", x"fa88", 
            x"ef5f", x"e2e1", x"e767", x"ebc8", 
            x"e7c3", x"dcae", x"d968", x"e94c", 
            x"fab1", x"08f2", x"20c6", x"2dbb", 
            x"10bb", x"e119", x"dcb5", x"0897", 
            x"2675", x"18df", x"07c0", x"0bb4", 
            x"1bd2", x"29f0", x"2c39", x"30eb", 
            x"375c", x"2c90", x"1653", x"05ab", 
            x"0237", x"116d", x"1d29", x"15df", 
            x"1bd0", x"2c23", x"1d4c", x"fbbf", 
            x"f4b0", x"0da6", x"1c94", x"0965", 
            x"f635", x"f985", x"0790", x"1c1a", 
            x"253f", x"0dd0", x"f99f", x"083d", 
            x"11fb", x"fee9", x"ed36", x"f8ad", 
            x"1c2e", x"2a26", x"0afe", x"ebf3", 
            x"f430", x"180f", x"3825", x"37e1", 
            x"0853", x"d503", x"e381", x"1c04", 
            x"2ba2", x"012f", x"d75a", x"dc27", 
            x"f3fa", x"f3fd", x"ed2a", x"f6c8", 
            x"01fe", x"0cd4", x"1555", x"fd3b", 
            x"d3da", x"d549", x"008f", x"18b3", 
            x"0841", x"fc17", x"0532", x"006f", 
            x"f0fd", x"faf5", x"0cfb", x"0ab5", 
            x"0007", x"fb46", x"021e", x"0df9", 
            x"0fac", x"12fa", x"185e", x"130b", 
            x"1315", x"1d19", x"1811", x"0322", 
            x"f806", x"f558", x"e690", x"e45f", 
            x"0796", x"1250", x"defc", x"c301", 
            x"efa8", x"1eee", x"1a2f", x"f06d", 
            x"cd68", x"d47c", x"f727", x"0eb0", 
            x"0e81", x"f9ec", x"e482", x"e223", 
            x"ed98", x"ec14", x"d98e", x"d312", 
            x"d956", x"df97", x"ee87", x"f76b", 
            x"e637", x"e1a9", x"0105", x"12df", 
            x"fc31", x"ea40", x"f5e5", x"0345", 
            x"068f", x"0973", x"0b01", x"ff08", 
            x"edef", x"ed12", x"fba0", x"04cd", 
            x"028f", x"0141", x"08a7", x"110b", 
            x"10a0", x"02b7", x"ec94", x"e143", 
            x"e4ad", x"e5ce", x"d82d", x"d52d", 
            x"f6cb", x"1475", x"04b4", x"e0d6", 
            x"d6d4", x"ee2c", x"0132", x"fa15", 
            x"ee3c", x"f0b0", x"fdac", x"0147", 
            x"f5ce", x"f30c", x"0346", x"09e6", 
            x"f967", x"f2d8", x"0645", x"1cf9", 
            x"2980", x"2aa3", x"2ad8", x"2c1a", 
            x"2349", x"1eeb", x"2924", x"2a13", 
            x"1345", x"07c3", x"1c91", x"22a7", 
            x"0557", x"f31a", x"01da", x"109f", 
            x"06e0", x"f80b", x"fd00", x"0645", 
            x"f66b", x"e39e", x"f27b", x"020a", 
            x"f5e8", x"eede", x"f8c7", x"03bf", 
            x"0be0", x"1517", x"1c20", x"1451", 
            x"0833", x"0620", x"06e9", x"0bfe", 
            x"1d6d", x"266d", x"1e67", x"12c4", 
            x"084c", x"0859", x"1163", x"0e72", 
            x"f7bd", x"e9fc", x"fd19", x"202b", 
            x"3075", x"2056", x"fe50", x"efcd", 
            x"0629", x"194b", x"0b08", x"ef73", 
            x"e3a7", x"f27d", x"05bc", x"04d0", 
            x"fe15", x"f59d", x"e9df", x"fa07", 
            x"1538", x"0d0d", x"f4f0", x"edf8", 
            x"f8cf", x"fc5a", x"eac3", x"de84", 
            x"e1e2", x"e395", x"e00a", x"e4a1", 
            x"eef2", x"f823", x"f890", x"f4a8", 
            x"fb1a", x"fe18", x"ef1e", x"e524", 
            x"f0a8", x"010a", x"070a", x"036d", 
            x"054d", x"1369", x"2183", x"1881", 
            x"f7d4", x"e8ad", x"fa2f", x"0280", 
            x"ff0b", x"0558", x"0b5e", x"0822", 
            x"fedd", x"fc9c", x"0026", x"faf9", 
            x"0362", x"2978", x"3312", x"1545", 
            x"13d3", x"3257", x"2e95", x"02d8", 
            x"e62e", x"e197", x"e5f5", x"f580", 
            x"0535", x"fbc5", x"ecc0", x"fb47", 
            x"04c6", x"f2b2", x"eb01", x"f07f", 
            x"f099", x"f6a7", x"fb27", x"f632", 
            x"f0a6", x"ebb0", x"f6d5", x"12ed", 
            x"160d", x"ff21", x"fb84", x"0501", 
            x"0410", x"0c29", x"1709", x"0677", 
            x"ecd6", x"f348", x"0f11", x"0df3", 
            x"f7c6", x"f741", x"ff28", x"f25d", 
            x"eff1", x"0605", x"0819", x"ec19", 
            x"d1cb", x"d217", x"e522", x"f3b7", 
            x"fe3d", x"02e3", x"f787", x"f52b", 
            x"0704", x"14ec", x"081d", x"edad", 
            x"ebb8", x"f48c", x"e8bb", x"e739", 
            x"07e3", x"1b68", x"0c37", x"0449", 
            x"123d", x"13e7", x"fe49", x"ff76", 
            x"2748", x"37bb", x"1863", x"f991", 
            x"f240", x"f612", x"f8f2", x"f355", 
            x"f2ee", x"06c6", x"10c6", x"f7ae", 
            x"d855", x"e186", x"0a7a", x"1b7f", 
            x"05ba", x"de58", x"c8af", x"d9ea", 
            x"fa8c", x"0760", x"03af", x"ff76", 
            x"fcc2", x"fabb", x"f848", x"f664", 
            x"fb03", x"0765", x"0c2e", x"ff09", 
            x"eeb1", x"f895", x"16bf", x"2d24", 
            x"29fb", x"1347", x"08da", x"1859", 
            x"2803", x"2034", x"14d3", x"1967", 
            x"1d20", x"1847", x"1708", x"1a5d", 
            x"1809", x"180d", x"2489", x"2736", 
            x"1674", x"0d16", x"1140", x"16ff", 
            x"1fd1", x"2f2b", x"2ef4", x"0c27", 
            x"f7a1", x"0ea5", x"2010", x"110e", 
            x"ffc3", x"f8b6", x"e94b", x"d9aa", 
            x"e17f", x"f1d7", x"e6fa", x"dce4", 
            x"fb24", x"1d44", x"0ef4", x"edf9", 
            x"f159", x"05c4", x"fd9d", x"f6cc", 
            x"14f6", x"271c", x"1973", x"110b", 
            x"1020", x"07eb", x"f987", x"f66d", 
            x"0823", x"0ca9", x"ff13", x"0270", 
            x"0e89", x"0fea", x"1445", x"2312", 
            x"291b", x"1056", x"f0ea", x"f7cf", 
            x"15cd", x"13f6", x"ecce", x"ce79", 
            x"dfb0", x"019e", x"0397", x"f3f6", 
            x"fab7", x"16ad", x"16d3", x"f173", 
            x"e096", x"f638", x"0e35", x"1a24", 
            x"14a6", x"0555", x"057c", x"1628", 
            x"2462", x"271e", x"21cb", x"143b", 
            x"f7e2", x"da71", x"e97e", x"2202", 
            x"2aa4", x"e9f2", x"bf8e", x"e588", 
            x"18fe", x"0aa8", x"de74", x"d9bb", 
            x"ed0b", x"e91f", x"cfd0", x"cda5", 
            x"eacf", x"f1f6", x"dc28", x"d229", 
            x"d4de", x"ca55", x"b7aa", x"c16f", 
            x"e8d5", x"0112", x"ee66", x"d47e", 
            x"e051", x"0307", x"10e7", x"054e", 
            x"fa94", x"048f", x"2380", x"3dfd", 
            x"2c24", x"f671", x"e060", x"fe58", 
            x"1265", x"0050", x"f5f5", x"0237", 
            x"0549", x"ec97", x"d996", x"ed57", 
            x"0b4a", x"0e16", x"eda0", x"ccf5", 
            x"ddd0", x"14e8", x"2c89", x"0ac4", 
            x"dbaf", x"dc3e", x"0cd9", x"13de", 
            x"e412", x"d04d", x"ecfe", x"1609", 
            x"28b5", x"1116", x"ec8b", x"d94d", 
            x"e7e4", x"10ce", x"13cd", x"e2ac", 
            x"d3bf", x"fb05", x"08c2", x"f4da"
        ),
        -- Block 5
        (
            x"f5fb", x"094a", x"0ad3", x"fab9", 
            x"eff5", x"ef7e", x"f60d", x"0225", 
            x"fffb", x"f058", x"eadd", x"e9f7", 
            x"dd35", x"d9a1", x"f95a", x"1f27", 
            x"10ed", x"eb06", x"f2e2", x"177f", 
            x"1fba", x"08bd", x"0741", x"1cf1", 
            x"1b0c", x"0686", x"0748", x"17ce", 
            x"0da0", x"000b", x"14bb", x"1fea", 
            x"0edf", x"0973", x"144e", x"21fd", 
            x"27fc", x"19bd", x"fbea", x"e8d0", 
            x"f463", x"0b61", x"115d", x"043c", 
            x"00c8", x"1596", x"22de", x"108e", 
            x"fe14", x"0419", x"0734", x"f63e", 
            x"ec67", x"f8b6", x"fba9", x"e7de", 
            x"e419", x"f949", x"ff28", x"effa", 
            x"e3e1", x"f43f", x"1ddb", x"2b5b", 
            x"1196", x"060c", x"0d10", x"0858", 
            x"034a", x"0397", x"f468", x"dcfb", 
            x"e610", x"0f39", x"2913", x"21ba", 
            x"10d9", x"0a34", x"09a0", x"0db5", 
            x"1356", x"0894", x"f20e", x"e831", 
            x"ee3f", x"f39d", x"f9b7", x"08b0", 
            x"15ad", x"ffdf", x"cef4", x"c373", 
            x"d984", x"d4ed", x"c1ae", x"d59e", 
            x"07be", x"17c6", x"f21c", x"d02d", 
            x"e7d1", x"1e26", x"30a6", x"0f63", 
            x"e676", x"e4dd", x"f280", x"e664", 
            x"d224", x"dd53", x"fa98", x"ff97", 
            x"f35a", x"f384", x"0416", x"18b3", 
            x"1f5f", x"056e", x"e443", x"f33b", 
            x"1b65", x"0e74", x"d665", x"d0df", 
            x"00a0", x"055f", x"db85", x"dead", 
            x"027b", x"ef96", x"c57a", x"d599", 
            x"02b2", x"fd20", x"d058", x"c439", 
            x"e731", x"01b1", x"f7ac", x"e75a", 
            x"e661", x"e217", x"de3f", x"f6ab", 
            x"1121", x"01b4", x"e8de", x"f719", 
            x"0fda", x"101d", x"fd77", x"f31a", 
            x"05ea", x"27f0", x"388d", x"255f", 
            x"07cb", x"0a65", x"1f73", x"2ef8", 
            x"40ea", x"39dc", x"1538", x"fa3f", 
            x"f048", x"f35c", x"0b1e", x"1f84", 
            x"083e", x"da7e", x"c9ec", x"dbd6", 
            x"f5de", x"fdd6", x"f13d", x"e7f6", 
            x"e040", x"d5fb", x"eb4d", x"0d3e", 
            x"fbba", x"d12a", x"d2fe", x"f6d2", 
            x"02a1", x"eaf9", x"d22a", x"dd6c", 
            x"03b1", x"0602", x"e0eb", x"d6a4", 
            x"f225", x"14a3", x"2a0f", x"2b36", 
            x"289a", x"29a5", x"2016", x"1986", 
            x"349f", x"4635", x"2728", x"0afa", 
            x"1f11", x"3eab", x"41f5", x"345e", 
            x"26a8", x"1cd9", x"1192", x"1a09", 
            x"2efb", x"225d", x"034a", x"10ae", 
            x"3f6b", x"498f", x"264f", x"0d58", 
            x"0216", x"e396", x"d4be", x"f1be", 
            x"0bcc", x"fc45", x"dfda", x"d483", 
            x"e682", x"0455", x"0b01", x"fd09", 
            x"e79a", x"d5de", x"d65a", x"efb0", 
            x"0967", x"05fc", x"f481", x"f697", 
            x"09bc", x"0eca", x"fd31", x"f7b2", 
            x"1271", x"24bc", x"171a", x"0d3b", 
            x"18fc", x"1b8e", x"0a3e", x"02d2", 
            x"0c7b", x"0402", x"ecab", x"f34e", 
            x"0ef8", x"113a", x"01dd", x"0b18", 
            x"2682", x"2f99", x"1b87", x"0924", 
            x"1871", x"3694", x"2ed2", x"0475", 
            x"ec7c", x"ff07", x"143c", x"f4ed", 
            x"c1f9", x"c417", x"eec4", x"f8de", 
            x"dd6f", x"d844", x"f24b", x"075b", 
            x"0948", x"ff25", x"f32a", x"f988", 
            x"1790", x"25d2", x"110f", x"fe28", 
            x"0a55", x"20a6", x"1e86", x"049e", 
            x"f2ff", x"03c4", x"1cef", x"1ef2", 
            x"0cc8", x"02e0", x"18b7", x"30e2", 
            x"2004", x"fc72", x"efee", x"f12c", 
            x"0074", x"1572", x"1a65", x"107e", 
            x"f6bb", x"e480", x"f955", x"0651", 
            x"f12b", x"e778", x"f918", x"0cb3", 
            x"0624", x"ed10", x"e2b4", x"f730", 
            x"0d25", x"1821", x"1b8d", x"0c24", 
            x"0242", x"0c4f", x"1a13", x"264c", 
            x"2f43", x"2eae", x"20b1", x"0b92", 
            x"030d", x"0e6b", x"136a", x"12a5", 
            x"1de6", x"1b06", x"fbb5", x"e55c", 
            x"f0f1", x"fede", x"f060", x"ebcf", 
            x"0c72", x"1a34", x"f4e1", x"da63", 
            x"e1bf", x"e029", x"e3b1", x"016c", 
            x"0f14", x"ef2a", x"c9a0", x"cbe5", 
            x"eb95", x"015d", x"ffe1", x"fb36", 
            x"067f", x"0f58", x"0132", x"f792", 
            x"00f3", x"129a", x"1855", x"f6f4", 
            x"c39b", x"be1b", x"e3e1", x"fad2", 
            x"f895", x"fa42", x"fd97", x"f5bd", 
            x"f0e1", x"005e", x"0bc7", x"f93f", 
            x"dd82", x"dd41", x"edef", x"e6b7", 
            x"cd95", x"d237", x"fba3", x"16a9", 
            x"0640", x"dd29", x"cd83", x"e75b", 
            x"f8c4", x"e800", x"de78", x"f3d1", 
            x"05e1", x"f989", x"e9d7", x"ef96", 
            x"f5b3", x"f2b0", x"fd06", x"0f12", 
            x"fbb3", x"d3f9", x"cf18", x"e6a1", 
            x"f118", x"e8ad", x"e182", x"e134", 
            x"e007", x"de96", x"e7f9", x"f856", 
            x"fd4d", x"f393", x"e9b0", x"dbfc", 
            x"d5f7", x"f096", x"fa68", x"d725", 
            x"ca3f", x"e381", x"f2b2", x"f506", 
            x"fdfb", x"ff4f", x"f27f", x"ece3", 
            x"f77f", x"ff21", x"f420", x"ef2b", 
            x"00e8", x"02b1", x"f115", x"ed3d", 
            x"0963", x"270a", x"1d21", x"033a", 
            x"ff20", x"0c24", x"1b50", x"2c0a", 
            x"30ce", x"2b0c", x"2575", x"11c0", 
            x"f27e", x"ef23", x"0c68", x"29f8", 
            x"234e", x"0c65", x"1bec", x"34c6", 
            x"285f", x"1736", x"1e01", x"1fbd", 
            x"0c85", x"fc8f", x"fa9a", x"f7c2", 
            x"0066", x"0fb2", x"0430", x"fe13", 
            x"1dbd", x"2ba7", x"0e63", x"f229", 
            x"f642", x"18c8", x"2a2b", x"0993", 
            x"ef50", x"fd4e", x"1121", x"29cb", 
            x"3ffb", x"2d69", x"1359", x"240b", 
            x"35df", x"20fb", x"fdf5", x"f9a9", 
            x"1c70", x"2aad", x"0d44", x"fda0", 
            x"0b5e", x"1862", x"1a22", x"0c67", 
            x"fc4c", x"0b17", x"19a4", x"0f89", 
            x"0bea", x"1733", x"2131", x"09b0", 
            x"ebb8", x"fed7", x"1e6b", x"1459", 
            x"fa50", x"f415", x"135d", x"302e", 
            x"11dd", x"f3e8", x"0919", x"17fb", 
            x"0c1d", x"045a", x"026f", x"03bb", 
            x"04f7", x"f9a3", x"e093", x"d13b", 
            x"de7e", x"ea94", x"e22e", x"dc1c", 
            x"e5f6", x"0166", x"1bfc", x"168e", 
            x"0455", x"0701", x"0f1e", x"12c7", 
            x"20cb", x"274d", x"0896", x"e0ad", 
            x"dc4e", x"fd94", x"0ce5", x"eaad", 
            x"c553", x"ce92", x"f229", x"fcb5", 
            x"e9d9", x"dfaa", x"f227", x"03e0", 
            x"fafe", x"ef85", x"f57b", x"fd5a", 
            x"fd8c", x"f323", x"def9", x"df3e", 
            x"048a", x"1ecc", x"09d8", x"e450", 
            x"de08", x"f0b8", x"e67d", x"cbf0", 
            x"d1b1", x"eb72", x"ee3a", x"e3d5", 
            x"e983", x"de4f", x"c299", x"c74b", 
            x"e6be", x"f4ff", x"eb3a", x"d242", 
            x"c9b3", x"e457", x"fc17", x"fc4e", 
            x"fe98", x"0d51", x"0f33", x"02a8", 
            x"f46f", x"eeb8", x"fc4a", x"165b", 
            x"234c", x"1e62", x"12fa", x"0993", 
            x"059c", x"025c", x"0178", x"05e0", 
            x"00cc", x"ea3c", x"ec2c", x"1881", 
            x"3643", x"2c3e", x"166d", x"fec5", 
            x"f760", x"0920", x"045c", x"ed02", 
            x"f121", x"fcae", x"f3be", x"e195", 
            x"dc4c", x"eac4", x"ef7c", x"d585", 
            x"d159", x"04cb", x"295b", x"1396", 
            x"f764", x"fcd9", x"055b", x"f321", 
            x"e44b", x"ee95", x"fece", x"fb51", 
            x"f5e4", x"0646", x"2466", x"38aa", 
            x"241a", x"02da", x"04c0", x"1bf5", 
            x"1d19", x"0ff8", x"0ccd", x"16aa", 
            x"24ad", x"1b3c", x"ff55", x"f83e", 
            x"012e", x"fb05", x"f5e1", x"f37b", 
            x"df7d", x"d790", x"ec19", x"01d5", 
            x"0536", x"fd36", x"f142", x"efec", 
            x"0f6a", x"3097", x"29f7", x"10ca", 
            x"fd20", x"e895", x"e3a3", x"f282", 
            x"e6ff", x"c50f", x"ba09", x"d4c0", 
            x"fe9e", x"08da", x"fe49", x"101a", 
            x"2726", x"06cf", x"dc38", x"f052", 
            x"1c22", x"1977", x"f676", x"e7d0", 
            x"f4d1", x"0a3b", x"1fa5", x"29c2", 
            x"1ee5", x"075a", x"fa3c", x"0c20", 
            x"1ca6", x"1770", x"0744", x"eb86", 
            x"e14a", x"0567", x"2107", x"12ce", 
            x"0806", x"0c0a", x"0e44", x"18b2", 
            x"2542", x"21e7", x"168d", x"08a8", 
            x"fe57", x"00e7", x"0e12", x"1b78", 
            x"1a28", x"14b5", x"2e2b", x"4180", 
            x"296f", x"147e", x"1b55", x"2706", 
            x"1c40", x"f84a", x"f2d3", x"102b", 
            x"09e3", x"ff4b", x"1e2d", x"1f1f", 
            x"f339", x"da58", x"dd2b", x"ebda", 
            x"ff36", x"09d1", x"0f2b", x"0c74", 
            x"1014", x"1b78", x"1426", x"01e4", 
            x"02be", x"1557", x"2355", x"1892", 
            x"0a21", x"1a09", x"1ae4", x"fc37", 
            x"ff40", x"29e3", x"351b", x"0df2", 
            x"f67e", x"0bb4", x"180c", x"2002", 
            x"3fb9", x"4859", x"2a84", x"0bfa", 
            x"04c9", x"0d9e", x"0ebc", x"fd33", 
            x"f380", x"0e33", x"1c35", x"fb0f", 
            x"d8e7", x"e180", x"039c", x"148d", 
            x"0459", x"db57", x"c215", x"d1b0", 
            x"f552", x"0a06", x"00dd", x"e546", 
            x"de8f", x"f835", x"0247", x"f9b9", 
            x"fb05", x"f990", x"014e", x"1acc", 
            x"1b15", x"0a33", x"13fb", x"2bdb", 
            x"2ca6", x"1fcd", x"19c9", x"20d9", 
            x"2bdd", x"2090", x"0d77", x"1062", 
            x"127b", x"fd74", x"f002", x"0102", 
            x"03a8", x"dfa0", x"d263", x"f49d", 
            x"08ed", x"ebed", x"c9b9", x"d47c", 
            x"e689", x"dca7", x"d337", x"e1b3", 
            x"f8ce", x"0319", x"051e", x"fc94", 
            x"e37a", x"d3bb", x"ec52", x"11da", 
            x"050d", x"c581", x"a731", x"cf51", 
            x"0176", x"0e05", x"063b", x"fd6a", 
            x"f739", x"ebdf", x"de48", x"e5dc", 
            x"fdd8", x"fd58", x"f75a", x"098f", 
            x"157f", x"0c8d", x"027a", x"fc1c", 
            x"f1cb", x"faf1", x"fbc0", x"e091", 
            x"dd0a", x"035e", x"2622", x"1dee", 
            x"f04f", x"d0b2", x"e4fa", x"0750", 
            x"03d3", x"de38", x"d528", x"0661", 
            x"30f0", x"1500", x"f0ee", x"1168", 
            x"47cc", x"42c7", x"fe6b", x"cfa6", 
            x"e5b0", x"ee82", x"c069", x"a244", 
            x"ceaa", x"0bda", x"0398", x"d9c8", 
            x"d6ef", x"ea06", x"e2e5", x"d727", 
            x"dff2", x"de57", x"cd0f", x"c40a", 
            x"c6ec", x"d678", x"f4ad", x"0a73", 
            x"f807", x"e11f", x"f7fe", x"2556", 
            x"308b", x"0b6c", x"f0e5", x"02fe", 
            x"0fb2", x"036e", x"008f", x"1570", 
            x"20bf", x"080b", x"f54a", x"0926", 
            x"21f5", x"1426", x"fb38", x"0566", 
            x"2205", x"16c3", x"f758", x"ffcf", 
            x"0db0", x"f5da", x"e2ec", x"e80e", 
            x"e0e1", x"c6fc", x"b9da", x"cf22", 
            x"f78b", x"08ac", x"ed96", x"dc62", 
            x"e724", x"de0f", x"cc30", x"d564", 
            x"e348", x"ef2d", x"00ea", x"f7fe", 
            x"f009", x"0b1a", x"2658", x"0f09", 
            x"dadf", x"dab0", x"153a", x"278c", 
            x"f8e1", x"e6f3", x"002c", x"0a64", 
            x"0fa5", x"1b98", x"13fc", x"ff27", 
            x"f6f3", x"0537", x"168f", x"0d9c", 
            x"f276", x"f69f", x"0a51", x"0938", 
            x"f95b", x"f383", x"ff1c", x"10b5", 
            x"14d4", x"ff2d", x"dba1", x"bc4e", 
            x"b837", x"d8b1", x"f7d2", x"0a07", 
            x"1156", x"fdea", x"004d", x"2603", 
            x"261b", x"040c", x"061c", x"1760", 
            x"0840", x"fb61", x"1414", x"361a", 
            x"2ac2", x"00b3", x"0276", x"29b5", 
            x"3041", x"159a", x"07af", x"06b8", 
            x"0ac6", x"1b82", x"272f", x"156e", 
            x"fd5d", x"fd53", x"0907", x"0a13", 
            x"fe17", x"ea75", x"d82f", x"daf1", 
            x"eaac", x"fce8", x"f850", x"d998", 
            x"efb4", x"2eea", x"3144", x"0a17", 
            x"088c", x"1d5b", x"1ecc", x"0e5e", 
            x"ff86", x"fd3c", x"0806", x"1f6e", 
            x"3426", x"2471", x"fd42", x"fbdd"
        ),
        -- Block 4
        (
            x"2175", x"3b78", x"3039", x"271d", 
            x"2bd0", x"0adb", x"e5d3", x"080d", 
            x"451d", x"4c08", x"209f", x"ef98", 
            x"d605", x"dd60", x"fc91", x"0e7a", 
            x"fa55", x"dfc3", x"d6ef", x"da75", 
            x"e113", x"f17f", x"016b", x"f151", 
            x"c8bf", x"bea0", x"e8b8", x"023a", 
            x"de30", x"cbd0", x"0034", x"1dc0", 
            x"f3ed", x"dd8b", x"077b", x"202e", 
            x"0035", x"f0d1", x"09ba", x"237b", 
            x"1e33", x"f7ea", x"e9ce", x"1535", 
            x"30fe", x"1579", x"fe6c", x"05fe", 
            x"0d15", x"0582", x"e970", x"d465", 
            x"eb1c", x"0020", x"ef47", x"db7b", 
            x"ecf5", x"1316", x"1651", x"f8d9", 
            x"e539", x"ecab", x"fc04", x"f942", 
            x"ee9d", x"f199", x"f916", x"eba6", 
            x"d2f9", x"d9f7", x"07af", x"21a5", 
            x"0995", x"ea0c", x"e8d6", x"0771", 
            x"2c32", x"27e7", x"fa73", x"ed89", 
            x"1065", x"1491", x"f387", x"e5a3", 
            x"01f4", x"2479", x"1067", x"ecfe", 
            x"fd3a", x"15cd", x"0bfb", x"0090", 
            x"fdaf", x"efee", x"e548", x"f706", 
            x"244e", x"244d", x"f67d", x"f5ac", 
            x"0816", x"ef15", x"d792", x"ef1a", 
            x"1225", x"110d", x"f258", x"e28f", 
            x"f52e", x"0b7d", x"0669", x"f4e4", 
            x"e9fd", x"e1dd", x"da61", x"e5fb", 
            x"0617", x"1818", x"0a72", x"e8bb", 
            x"ddee", x"025b", x"21af", x"124d", 
            x"f9e5", x"012f", x"2594", x"4193", 
            x"2d6d", x"01f9", x"fb36", x"1ed7", 
            x"380c", x"262e", x"0960", x"fec7", 
            x"0c3b", x"270d", x"3c21", x"3a20", 
            x"241c", x"0ee9", x"ef81", x"e306", 
            x"011b", x"1479", x"ffc1", x"ef0c", 
            x"e492", x"cf65", x"da0c", x"0d9a", 
            x"30b1", x"261a", x"01f3", x"ea86", 
            x"fd2b", x"1489", x"ffe5", x"e972", 
            x"ffe5", x"06a4", x"ed36", x"eeac", 
            x"ff16", x"ff02", x"009a", x"0a63", 
            x"0f18", x"15aa", x"0e76", x"004f", 
            x"03c1", x"10b3", x"11f3", x"f631", 
            x"eafa", x"1297", x"31dc", x"18ab", 
            x"e7e4", x"d94f", x"ff25", x"213f", 
            x"1652", x"0939", x"0001", x"f252", 
            x"017a", x"20a1", x"11f4", x"dc69", 
            x"cd21", x"f275", x"1913", x"2a81", 
            x"2288", x"fd31", x"e603", x"018a", 
            x"2639", x"176f", x"f70b", x"f840", 
            x"00d5", x"f84f", x"099d", x"25bc", 
            x"11ec", x"ef78", x"f77f", x"069d", 
            x"f07f", x"e09a", x"ee33", x"f75d", 
            x"ea59", x"df82", x"e8eb", x"fd6e", 
            x"0643", x"03cc", x"f176", x"cd67", 
            x"be5a", x"e04d", x"f62a", x"d71a", 
            x"c2f6", x"e6b4", x"10e8", x"1323", 
            x"026b", x"00c0", x"0b96", x"05e7", 
            x"dd61", x"bde7", x"c5aa", x"c5d8", 
            x"b9dc", x"d48e", x"fd43", x"f973", 
            x"dd55", x"e8f3", x"1638", x"2122", 
            x"feef", x"eb0b", x"eb6f", x"e845", 
            x"0157", x"2401", x"20ec", x"08fc", 
            x"00e4", x"0f91", x"2655", x"1d7b", 
            x"0184", x"006e", x"07b3", x"f91a", 
            x"ef7f", x"f3cc", x"fc22", x"109d", 
            x"1764", x"0a29", x"fc11", x"f064", 
            x"f0f5", x"0546", x"12bc", x"fe36", 
            x"e5c8", x"f3ec", x"0bd9", x"fc40", 
            x"e713", x"f60d", x"0c0d", x"fdc2", 
            x"d633", x"c9aa", x"f666", x"18aa", 
            x"f9ec", x"f158", x"135c", x"157e", 
            x"f4c7", x"df99", x"f110", x"1cab", 
            x"2dd4", x"1578", x"01f8", x"192c", 
            x"3022", x"1921", x"fbcf", x"05ee", 
            x"28cc", x"346b", x"15cf", x"f66e", 
            x"1261", x"3c4a", x"2609", x"f91b", 
            x"f9fa", x"14dd", x"23b4", x"2298", 
            x"228b", x"0e42", x"f80d", x"0362", 
            x"0edc", x"0caa", x"12d8", x"0c2c", 
            x"ea65", x"e3fe", x"1856", x"4146", 
            x"11c4", x"dbaa", x"f70b", x"315f", 
            x"31b1", x"fadf", x"f011", x"2d6c", 
            x"4df2", x"2162", x"ef83", x"ff4d", 
            x"23f8", x"0575", x"ce70", x"dde2", 
            x"17fc", x"28f6", x"13a9", x"0198", 
            x"020f", x"0c2f", x"1b40", x"21a4", 
            x"0fce", x"f652", x"ed56", x"f9f0", 
            x"0596", x"f906", x"de7e", x"e16a", 
            x"f9ea", x"fb32", x"e104", x"e340", 
            x"ff72", x"0640", x"fd69", x"f22c", 
            x"eaff", x"f58c", x"19cc", x"2728", 
            x"104f", x"0d53", x"1ee4", x"3594", 
            x"3947", x"0b58", x"ed3e", x"10e9", 
            x"38c7", x"3226", x"0ee4", x"faa8", 
            x"0875", x"1abd", x"19c4", x"06d9", 
            x"fb20", x"0a84", x"158c", x"fed7", 
            x"fc15", x"10ab", x"08d8", x"f833", 
            x"0342", x"2809", x"1ddd", x"ec8d", 
            x"ee50", x"1832", x"14e3", x"f651", 
            x"fbbd", x"14bb", x"106a", x"06bd", 
            x"223c", x"313e", x"0ce6", x"f87b", 
            x"0bf9", x"fc1a", x"d86a", x"dfad", 
            x"f42d", x"f08f", x"ef2c", x"f859", 
            x"0e0a", x"1742", x"097c", x"0815", 
            x"0d32", x"0e84", x"20e0", x"2825", 
            x"056d", x"e04d", x"f291", x"1d92", 
            x"1721", x"fde9", x"023a", x"00fa", 
            x"eb17", x"ec95", x"002f", x"f33f", 
            x"db94", x"e7c6", x"e6f2", x"c61d", 
            x"d43e", x"145f", x"363a", x"0c48", 
            x"d519", x"d590", x"e2fd", x"db2b", 
            x"e58f", x"012f", x"f9b1", x"d131", 
            x"bdf3", x"dd15", x"0b56", x"ff2e", 
            x"d1c6", x"d580", x"ef90", x"ed74", 
            x"eee2", x"ff69", x"fbf3", x"ee40", 
            x"f403", x"0a04", x"1668", x"f823", 
            x"d529", x"da43", x"f847", x"0795", 
            x"ee88", x"dbb4", x"e14f", x"e653", 
            x"f385", x"06ab", x"0153", x"f1c8", 
            x"feec", x"0e8a", x"042a", x"f2bb", 
            x"ed8f", x"e81b", x"dd5b", x"dfca", 
            x"f128", x"f65c", x"ed25", x"f64f", 
            x"06d8", x"0ff0", x"19de", x"1df4", 
            x"03cd", x"ee41", x"078d", x"206d", 
            x"f99b", x"bd3f", x"b5fc", x"d453", 
            x"eccf", x"e724", x"ea47", x"0c7a", 
            x"fc43", x"aea3", x"915f", x"c031", 
            x"ec7a", x"e79e", x"c714", x"afab", 
            x"b6a4", x"c3d0", x"df6d", x"1107", 
            x"1bc4", x"f223", x"c955", x"cf8d", 
            x"f2d0", x"f67e", x"e969", x"fe67", 
            x"0d24", x"08d0", x"0a63", x"097f", 
            x"0a8b", x"145d", x"169e", x"184b", 
            x"0e6c", x"fca6", x"ff61", x"0caf", 
            x"1273", x"1162", x"0c0a", x"08e7", 
            x"1d80", x"2bec", x"0e20", x"ecac", 
            x"001e", x"378f", x"516c", x"26f4", 
            x"e9f1", x"efa3", x"2a1a", x"47b1", 
            x"1749", x"db24", x"da99", x"094a", 
            x"216d", x"fdce", x"e70f", x"0014", 
            x"1409", x"075f", x"fbd4", x"05c1", 
            x"1145", x"21ef", x"3415", x"1b25", 
            x"e839", x"e507", x"2366", x"41fd", 
            x"f86c", x"b109", x"d7e1", x"2617", 
            x"2886", x"02b3", x"072c", x"134c", 
            x"fcce", x"edcd", x"f5a8", x"0052", 
            x"fda2", x"db92", x"c122", x"e328", 
            x"0fcd", x"0a4e", x"ee65", x"eaa4", 
            x"06a4", x"1a57", x"f9c8", x"d3f7", 
            x"f727", x"1919", x"03cd", x"f37b", 
            x"02b2", x"0b87", x"0738", x"17a2", 
            x"28de", x"2516", x"220a", x"1cab", 
            x"0658", x"0f35", x"1ec6", x"10b9", 
            x"0712", x"0137", x"feea", x"094f", 
            x"1b47", x"1d18", x"121c", x"ff4b", 
            x"f8f2", x"034c", x"1582", x"30b8", 
            x"3447", x"1d33", x"02fb", x"ee74", 
            x"fe7f", x"293a", x"2d58", x"0885", 
            x"e217", x"ed62", x"2e1a", x"4fab", 
            x"2923", x"f28d", x"de3c", x"eeed", 
            x"054f", x"08c9", x"f6ba", x"eab6", 
            x"ecb7", x"00d2", x"14bf", x"1559", 
            x"0a8e", x"ecea", x"ea43", x"0e50", 
            x"056c", x"d89e", x"e417", x"21aa", 
            x"390d", x"fb1e", x"c689", x"e9f9", 
            x"0c40", x"dd67", x"b885", x"e588", 
            x"0c79", x"f7fc", x"db0e", x"dade", 
            x"e576", x"e9ba", x"e4ca", x"e3ad", 
            x"ec22", x"e922", x"e160", x"ebcd", 
            x"01fd", x"0eb6", x"0948", x"f3db", 
            x"e69a", x"07d2", x"24fc", x"0114", 
            x"e388", x"0443", x"33a4", x"331d", 
            x"0ba4", x"f8e0", x"f738", x"e820", 
            x"e679", x"fe73", x"1d24", x"16be", 
            x"e625", x"e06b", x"1a80", x"2ebb", 
            x"f9a2", x"dcca", x"f8d3", x"0d66", 
            x"00fc", x"f58c", x"0ba7", x"2753", 
            x"1221", x"db2f", x"d9f9", x"196f", 
            x"3314", x"fee7", x"cfb3", x"d78c", 
            x"fce7", x"1727", x"fbe4", x"e786", 
            x"0cbc", x"1710", x"f0f2", x"e60b", 
            x"f741", x"0353", x"07e1", x"0451", 
            x"ed6e", x"dc9e", x"f5bd", x"0c2f", 
            x"ec18", x"d431", x"eb2b", x"03d8", 
            x"176b", x"1eca", x"0d17", x"f5e5", 
            x"de1d", x"e77b", x"19c5", x"215d", 
            x"f814", x"f03a", x"1354", x"25a0", 
            x"1577", x"0dd2", x"11c4", x"02fc", 
            x"e94c", x"ee55", x"0284", x"fb3b", 
            x"f464", x"0724", x"1f22", x"139f", 
            x"01cc", x"19b3", x"291d", x"0b24", 
            x"fb63", x"021b", x"06fe", x"1510", 
            x"2075", x"0cb6", x"ec45", x"e2da", 
            x"f9e1", x"0c06", x"fc20", x"f5cf", 
            x"0e2b", x"1368", x"f52c", x"e709", 
            x"ff5f", x"1cc1", x"14ba", x"fd52", 
            x"0718", x"16a4", x"0d06", x"0635", 
            x"0a9e", x"0d79", x"09d6", x"f150", 
            x"d654", x"e6fc", x"1ba5", x"3698", 
            x"0c2d", x"e71f", x"178b", x"3d4a", 
            x"0a9a", x"e64c", x"0462", x"17ae", 
            x"0ed5", x"1116", x"277f", x"300f", 
            x"1172", x"ebc1", x"f24a", x"0339", 
            x"f466", x"e8a8", x"fcd5", x"124d", 
            x"1663", x"1f9e", x"155d", x"fa7b", 
            x"f4ca", x"fe22", x"f454", x"ee79", 
            x"fd15", x"036a", x"0413", x"fa90", 
            x"0c5a", x"286a", x"1c73", x"ff37", 
            x"fea2", x"0fc3", x"ff5f", x"dc82", 
            x"e3d9", x"fb06", x"fe89", x"fd68", 
            x"f6fc", x"e8bc", x"ea37", x"025f", 
            x"0894", x"ecab", x"de8a", x"eb77", 
            x"f700", x"f4c4", x"e23a", x"bda6", 
            x"b84e", x"e5aa", x"04c0", x"ddee", 
            x"ae8b", x"cc7d", x"fa25", x"fcce", 
            x"fa93", x"fafd", x"f118", x"fccf", 
            x"0e25", x"fe15", x"e912", x"ec28", 
            x"0597", x"19ec", x"139a", x"0c56", 
            x"1234", x"1d08", x"24bb", x"3155", 
            x"393f", x"278b", x"fac1", x"dd68", 
            x"f750", x"25a7", x"18d4", x"f21f", 
            x"0275", x"1953", x"0837", x"fb33", 
            x"fe91", x"e5d1", x"c806", x"dc59", 
            x"12e0", x"226c", x"f7da", x"dc3d", 
            x"e4d4", x"e088", x"cde8", x"dc62", 
            x"facf", x"fae1", x"e23d", x"d1b9", 
            x"e9aa", x"0dcb", x"07bd", x"f3d9", 
            x"f00b", x"ea30", x"e50b", x"cadc", 
            x"b915", x"ee2a", x"20ce", x"f6b6", 
            x"b33e", x"adf4", x"d493", x"f842", 
            x"fa77", x"e969", x"cbcb", x"b3c3", 
            x"cea4", x"fa79", x"f168", x"d0f1", 
            x"d4b1", x"f42a", x"0659", x"f17c", 
            x"ddb3", x"e3a6", x"e630", x"f47a", 
            x"1522", x"0cde", x"e814", x"e79a", 
            x"fcd2", x"1f89", x"3f57", x"4be8", 
            x"3473", x"0a49", x"10b3", x"483c", 
            x"5f71", x"4b6b", x"3000", x"2166", 
            x"3870", x"4e04", x"3cb8", x"16d7", 
            x"144a", x"2df4", x"4318", x"3e53", 
            x"2209", x"189b", x"1d6d", x"0aab", 
            x"fdce", x"2bdc", x"3d5a", x"f8e2", 
            x"c26d", x"d66d", x"0021", x"0cc1", 
            x"03d6", x"f956", x"ffd9", x"06f5", 
            x"02ee", x"0474", x"fb97", x"f511", 
            x"090e", x"1506", x"0722", x"0246", 
            x"0534", x"f4f8", x"f1a7", x"154f", 
            x"41f2", x"3d1a", x"0f59", x"1685", 
            x"38d6", x"294d", x"259b", x"49bb", 
            x"3c9a", x"fb32", x"d439", x"e451", 
            x"f5bd", x"eb6c", x"07a9", x"3662", 
            x"13d1", x"d176", x"d64c", x"ffe2", 
            x"ffe0", x"dcb3", x"deb4", x"18ae", 
            x"254c", x"d71c", x"a8dd", x"ec57"
        ),
        -- Block 3
        (
            x"35f6", x"2421", x"f87f", x"eb85", 
            x"e79e", x"f0d3", x"f6ec", x"ea13", 
            x"e362", x"e75c", x"f5ec", x"04d7", 
            x"f3e3", x"e61c", x"060c", x"2b93", 
            x"3005", x"2615", x"16d8", x"04ba", 
            x"012d", x"1b6c", x"2d65", x"10c5", 
            x"03b6", x"2e74", x"4a31", x"23a7", 
            x"f979", x"15a1", x"4bce", x"26cd", 
            x"d48b", x"d56d", x"12f2", x"2dca", 
            x"2518", x"17e5", x"fab7", x"e65d", 
            x"f1c8", x"f71e", x"e7b5", x"db5e", 
            x"d8b3", x"d02b", x"cccd", x"d4f4", 
            x"d147", x"e18b", x"0b1e", x"12d3", 
            x"df2d", x"b7ff", x"d6db", x"fc71", 
            x"ee9c", x"cf0f", x"db0b", x"f680", 
            x"e9ca", x"d5ed", x"d9a5", x"ed76", 
            x"095b", x"1a43", x"10f2", x"0630", 
            x"fc09", x"efbf", x"ef87", x"fa89", 
            x"0a55", x"25c3", x"3ee0", x"35a5", 
            x"28da", x"2ea1", x"31aa", x"3a5d", 
            x"4687", x"2dcc", x"0dea", x"07ab", 
            x"10f2", x"1577", x"13fd", x"2724", 
            x"3ac5", x"1eb5", x"0154", x"106c", 
            x"2452", x"2841", x"150d", x"086c", 
            x"0903", x"f813", x"e4f0", x"e328", 
            x"ee4e", x"00a7", x"1642", x"0d8d", 
            x"ebd7", x"ee31", x"18ff", x"37df", 
            x"137c", x"d80c", x"d977", x"013e", 
            x"f430", x"ce28", x"e74b", x"0faf", 
            x"fe1c", x"d9a4", x"d4ea", x"ef6c", 
            x"1176", x"0808", x"e2f4", x"e54b", 
            x"10b7", x"34f2", x"259a", x"e123", 
            x"c582", x"fc88", x"27e1", x"1233", 
            x"f1b0", x"f967", x"0d5b", x"0849", 
            x"f399", x"dc93", x"e71b", x"2263", 
            x"249d", x"d0fa", x"ab3e", x"db95", 
            x"01b1", x"f0e3", x"e7e8", x"0f27", 
            x"30d2", x"fce8", x"c8f0", x"f6de", 
            x"2f0e", x"1c99", x"f80e", x"03c0", 
            x"0f8b", x"11b5", x"0fa7", x"ee2e", 
            x"e5a5", x"2b28", x"4aa7", x"0b85", 
            x"cb34", x"cb2b", x"e879", x"e10b", 
            x"c1f7", x"e2cc", x"2339", x"08db", 
            x"c7c1", x"bc1b", x"cd21", x"cf1b", 
            x"d1c8", x"e107", x"d97b", x"c3cd", 
            x"d7d5", x"f4a9", x"f087", x"f6b2", 
            x"0dc3", x"0ca7", x"ffe4", x"0259", 
            x"fba4", x"ecc7", x"f6e4", x"177f", 
            x"2123", x"f783", x"d44e", x"f026", 
            x"0917", x"e519", x"d1d0", x"029a", 
            x"1da9", x"efe9", x"dfca", x"115a", 
            x"2a57", x"0055", x"d099", x"dce3", 
            x"0559", x"fc31", x"d13b", x"d989", 
            x"0866", x"047f", x"e7a6", x"f7f5", 
            x"050c", x"ee21", x"d5a4", x"ed63", 
            x"2100", x"2500", x"0461", x"f8bf", 
            x"0452", x"159f", x"1c83", x"162c", 
            x"106b", x"049c", x"02fa", x"0120", 
            x"ebf1", x"e39f", x"fb39", x"fc67", 
            x"d430", x"b4b4", x"ce15", x"1708", 
            x"1dd5", x"c97d", x"abf8", x"e922", 
            x"0759", x"fd85", x"f431", x"f768", 
            x"0936", x"05d6", x"03a0", x"266d", 
            x"266a", x"f26f", x"e91d", x"09ce", 
            x"065f", x"e1f7", x"dde9", x"0af5", 
            x"1c7b", x"04bf", x"02b3", x"132f", 
            x"1578", x"01af", x"f65f", x"215e", 
            x"503b", x"3ebc", x"0993", x"f999", 
            x"1932", x"32e6", x"2aca", x"1057", 
            x"0249", x"034d", x"137a", x"2527", 
            x"13d0", x"098f", x"0dc7", x"f6fc", 
            x"fba2", x"1ce1", x"0b0e", x"f684", 
            x"1124", x"1e9c", x"11bd", x"051d", 
            x"0217", x"0ea7", x"17fc", x"0b07", 
            x"f965", x"ffbd", x"09e7", x"03a1", 
            x"0777", x"11f9", x"fb1a", x"e01e", 
            x"f3dc", x"0324", x"e916", x"d54f", 
            x"dc7b", x"ec9b", x"f75b", x"f1a4", 
            x"ecd8", x"e426", x"d173", x"cae1", 
            x"00fe", x"2a69", x"e7f0", x"a136", 
            x"c832", x"19d5", x"197e", x"e7ac", 
            x"de04", x"fd67", x"fcad", x"e346", 
            x"e7fd", x"1aa3", x"3778", x"24da", 
            x"16a1", x"1c9f", x"1dec", x"1eee", 
            x"314a", x"3456", x"13c2", x"0201", 
            x"2111", x"4988", x"3729", x"fa84", 
            x"f467", x"2e86", x"4e98", x"3039", 
            x"0f78", x"13a0", x"1f18", x"0a8d", 
            x"01ed", x"0c1d", x"fe1b", x"d115", 
            x"bccf", x"da5f", x"f781", x"e20e", 
            x"d474", x"f48b", x"f79a", x"ee35", 
            x"039d", x"fe66", x"d687", x"d818", 
            x"f51d", x"0f09", x"0f8f", x"ef1d", 
            x"f072", x"1c2f", x"2766", x"0ce2", 
            x"0977", x"1dae", x"2f8d", x"1902", 
            x"f14c", x"fa8f", x"2343", x"3aa6", 
            x"27f0", x"e339", x"b9c4", x"ea44", 
            x"1065", x"0216", x"f0d6", x"ea7f", 
            x"ee1a", x"fa76", x"ef68", x"dc43", 
            x"e3f4", x"fdd4", x"0b00", x"f98c", 
            x"e4a6", x"ebde", x"ff32", x"022c", 
            x"043a", x"f05c", x"dc15", x"e9c1", 
            x"024e", x"0e4e", x"fdd6", x"dfb2", 
            x"000b", x"4834", x"3fa7", x"067f", 
            x"13f0", x"372e", x"1949", x"fca7", 
            x"1824", x"42de", x"34b1", x"fa3d", 
            x"fb87", x"1e40", x"08ea", x"e53d", 
            x"fe9c", x"2471", x"14c9", x"eea5", 
            x"f83a", x"0949", x"de68", x"be01", 
            x"f2db", x"2ae5", x"fdf3", x"b9c6", 
            x"c7f2", x"eca2", x"e87b", x"d814", 
            x"cfbf", x"d21e", x"e126", x"f3b6", 
            x"f77d", x"f69f", x"f0e5", x"f93b", 
            x"09eb", x"0825", x"f332", x"fa7c", 
            x"18f7", x"13ba", x"09af", x"0f77", 
            x"2062", x"2d3f", x"1157", x"eb54", 
            x"f33a", x"2312", x"2eb9", x"028f", 
            x"d90e", x"e7b5", x"1280", x"109b", 
            x"f06f", x"d5dc", x"d724", x"f0f0", 
            x"fed7", x"f1bb", x"e1dd", x"f3d8", 
            x"1fea", x"1b21", x"e44f", x"cca1", 
            x"e5c2", x"0613", x"14cd", x"024d", 
            x"ddbc", x"cd5e", x"eef7", x"2406", 
            x"212e", x"ff09", x"f6ad", x"14c4", 
            x"3671", x"22be", x"f82f", x"ff12", 
            x"244a", x"2b25", x"0dfb", x"e1f5", 
            x"e1a4", x"0c34", x"1fe7", x"ffaf", 
            x"ef64", x"0b5b", x"021a", x"e141", 
            x"f0c3", x"0f60", x"eb76", x"ae45", 
            x"b107", x"d384", x"d8e7", x"e3fe", 
            x"0c8f", x"0fe3", x"d8a0", x"ca32", 
            x"094d", x"2a92", x"f5ec", x"d619", 
            x"e85e", x"feea", x"ff68", x"eec1", 
            x"fbad", x"0b75", x"0c0b", x"16d2", 
            x"2d94", x"1dab", x"09dd", x"0c57", 
            x"0968", x"0c3f", x"240c", x"3500", 
            x"285c", x"17c8", x"2540", x"41f4", 
            x"33aa", x"fea3", x"e350", x"e4e1", 
            x"dee2", x"e5ec", x"f51f", x"f4f3", 
            x"f5d9", x"e7da", x"d153", x"d791", 
            x"e248", x"e406", x"e50c", x"d9f7", 
            x"c772", x"dec0", x"0d13", x"1594", 
            x"eed8", x"d805", x"e928", x"fe14", 
            x"e3b4", x"c765", x"e502", x"fcc6", 
            x"f496", x"f65d", x"0b95", x"19ba", 
            x"0fd8", x"01d7", x"076e", x"199f", 
            x"2dae", x"286d", x"10dc", x"0adb", 
            x"1b06", x"3de3", x"54dc", x"3b3e", 
            x"17c2", x"10f0", x"247f", x"3669", 
            x"28de", x"0d45", x"1995", x"3e64", 
            x"303a", x"febe", x"fe40", x"379e", 
            x"49b2", x"0d52", x"dfd9", x"0cbd", 
            x"4bf5", x"2541", x"cdb9", x"d8d5", 
            x"218b", x"2784", x"ff40", x"fc23", 
            x"0d9f", x"fe74", x"ec74", x"10fc", 
            x"43a1", x"29d4", x"e5c2", x"e86a", 
            x"0ce0", x"0bc0", x"0a76", x"0af7", 
            x"f8d5", x"e89b", x"e87a", x"058d", 
            x"3272", x"37d3", x"177d", x"0eac", 
            x"2295", x"0381", x"d84e", x"f260", 
            x"23f3", x"2552", x"f406", x"beae", 
            x"c15f", x"f81e", x"0f09", x"f89c", 
            x"fecc", x"1aa9", x"145a", x"f22c", 
            x"d4e5", x"ea3b", x"28e7", x"2648", 
            x"f0bf", x"e3ea", x"f058", x"fefb", 
            x"03da", x"0ef4", x"2427", x"1581", 
            x"d9ae", x"c29f", x"f75a", x"2473", 
            x"09f7", x"dd95", x"e3da", x"f1f1", 
            x"0f30", x"36fe", x"1082", x"c8d1", 
            x"d828", x"0d9b", x"14c5", x"efa0", 
            x"d24b", x"ee06", x"12d9", x"14f3", 
            x"155a", x"09e4", x"f916", x"0754", 
            x"24c4", x"309b", x"1611", x"eaed", 
            x"ecc3", x"2194", x"1d99", x"f5ae", 
            x"ecdd", x"ec67", x"e25d", x"e63a", 
            x"dd59", x"bc9b", x"d1e5", x"1a16", 
            x"1503", x"c484", x"c589", x"16ed", 
            x"235a", x"f369", x"f8c7", x"1ba5", 
            x"1e89", x"f8f7", x"d066", x"dafb", 
            x"f10a", x"d87b", x"d8f3", x"f95b", 
            x"ef2b", x"e238", x"fb45", x"fdb0", 
            x"f714", x"027a", x"e64c", x"c565", 
            x"c977", x"caf0", x"ce0f", x"e924", 
            x"055d", x"ff7c", x"e30a", x"d3c6", 
            x"d777", x"ec63", x"ef16", x"c46e", 
            x"b2eb", x"cf91", x"e6ac", x"e9a1", 
            x"eb40", x"eb60", x"fcbc", x"07d0", 
            x"0483", x"0194", x"e1b2", x"ce35", 
            x"f22e", x"115c", x"18be", x"20ba", 
            x"0976", x"de32", x"f883", x"3ac2", 
            x"3461", x"faaf", x"de67", x"f7c4", 
            x"2212", x"2a75", x"10bf", x"0d20", 
            x"1dc9", x"1061", x"effa", x"e58a", 
            x"f9e9", x"1107", x"25af", x"3016", 
            x"25ec", x"0ff5", x"10d5", x"2169", 
            x"23e8", x"226d", x"1f66", x"253b", 
            x"35f7", x"3779", x"2701", x"2ade", 
            x"282b", x"1eb9", x"1d9f", x"11c8", 
            x"17d9", x"1f9b", x"e693", x"a91d", 
            x"be5a", x"faa9", x"0cac", x"d596", 
            x"a6cd", x"db81", x"244e", x"1fdf", 
            x"f0b9", x"c86b", x"cae4", x"127e", 
            x"307d", x"fd1f", x"d9c8", x"e6df", 
            x"12f1", x"3483", x"17ab", x"f397", 
            x"1391", x"39b9", x"3540", x"2442", 
            x"1147", x"fa0b", x"ef60", x"0740", 
            x"2467", x"fd55", x"c9c3", x"fc3f", 
            x"3642", x"1e5d", x"03d3", x"04a5", 
            x"15dd", x"156f", x"ee2b", x"e150", 
            x"fd8f", x"fd20", x"e2df", x"e111", 
            x"dfad", x"deb2", x"fd7a", x"22d5", 
            x"29bb", x"11cf", x"fe85", x"f933", 
            x"f88f", x"108f", x"2f15", x"0dd9", 
            x"f80d", x"30cf", x"43ff", x"03ad", 
            x"e01e", x"1d46", x"5ea4", x"463f", 
            x"0964", x"ed7b", x"027f", x"2e35", 
            x"3749", x"172e", x"ec94", x"e9a4", 
            x"1985", x"3adf", x"2374", x"f135", 
            x"d99f", x"e6f8", x"0e10", x"25b0", 
            x"16b5", x"f630", x"ec3a", x"f849", 
            x"fcc9", x"04bb", x"0932", x"f1b2", 
            x"d40b", x"e246", x"1594", x"1ae0", 
            x"f190", x"ed20", x"085b", x"0771", 
            x"dfe2", x"db2c", x"faf9", x"0ebe", 
            x"0c67", x"fdbb", x"f3a7", x"ec79", 
            x"0365", x"2757", x"0496", x"cc17", 
            x"dd49", x"1df4", x"218b", x"f7a4", 
            x"f0f7", x"10cc", x"0b1d", x"edcd", 
            x"0985", x"1f16", x"ee0c", x"c31f", 
            x"e3a3", x"0fd2", x"03d3", x"f950", 
            x"12bc", x"0c0e", x"d84c", x"abe4", 
            x"bfbd", x"edf4", x"e8a5", x"cfa9", 
            x"c5af", x"cc4f", x"dffc", x"e37f", 
            x"c5de", x"bcf6", x"e0b0", x"068c", 
            x"e8e7", x"b074", x"b438", x"f0b3", 
            x"2a48", x"2077", x"ee37", x"d528", 
            x"df99", x"f050", x"038e", x"00bf", 
            x"f9b3", x"085e", x"121d", x"0a66", 
            x"1874", x"1d7e", x"edee", x"d1e3", 
            x"f940", x"04e1", x"d7ea", x"c2f2", 
            x"f124", x"14c6", x"e6dc", x"b9bb", 
            x"ca56", x"ed13", x"007a", x"165e", 
            x"1025", x"d44d", x"b461", x"fa11", 
            x"4224", x"1b7a", x"e97f", x"0dc6", 
            x"1e41", x"df7c", x"c069", x"f836", 
            x"2948", x"2339", x"0d66", x"141e", 
            x"0b60", x"019e", x"3e6c", x"5595", 
            x"0eae", x"dce4", x"00ec", x"16cd", 
            x"ee53", x"db7b", x"01b2", x"2432", 
            x"0f2f", x"f93a", x"04d9", x"00e7", 
            x"02b1", x"0f00", x"f2ac", x"dc30", 
            x"0a81", x"2cc1", x"02d8", x"c0a1", 
            x"d400", x"0f32", x"00ed", x"ebad", 
            x"1bfe", x"3969", x"0f1e", x"f58e", 
            x"1e49", x"48c6", x"2e28", x"ff42", 
            x"0927", x"36eb", x"417d", x"2c20"
        ),
        -- Block 2
        (
            x"19e1", x"2174", x"32ec", x"2acc", 
            x"29a8", x"3a62", x"2b6b", x"0d27", 
            x"0424", x"0d85", x"1b20", x"1172", 
            x"00a2", x"07b2", x"2f71", x"41f2", 
            x"1ec8", x"fad8", x"fb37", x"0e19", 
            x"15b8", x"0461", x"f380", x"ff88", 
            x"f6bc", x"f9a7", x"1615", x"1f04", 
            x"1713", x"0100", x"ea88", x"f5c1", 
            x"054b", x"f6ae", x"ea23", x"eea6", 
            x"0c11", x"2e29", x"2166", x"ec19", 
            x"e588", x"0309", x"1a5a", x"182e", 
            x"fd87", x"fb38", x"1bd0", x"2469", 
            x"0116", x"16df", x"4798", x"1cba", 
            x"d8bc", x"fd7c", x"3e6a", x"0979", 
            x"a994", x"bd95", x"1842", x"2721", 
            x"eb5d", x"cc34", x"f175", x"18ce", 
            x"0f72", x"e9f3", x"dfc3", x"e10d", 
            x"c06b", x"c57f", x"f665", x"fa87", 
            x"dae8", x"d1e8", x"d313", x"dca8", 
            x"f2e0", x"0255", x"f651", x"c378", 
            x"c49d", x"11c8", x"2eaa", x"f501", 
            x"cfc3", x"e934", x"18f9", x"2759", 
            x"069e", x"059a", x"31f6", x"1e7b", 
            x"db4d", x"cbcb", x"ed86", x"0864", 
            x"fc72", x"e799", x"e41c", x"f226", 
            x"0657", x"fa78", x"e23f", x"e8bc", 
            x"edc0", x"dbbc", x"d857", x"e220", 
            x"e94a", x"0105", x"0bdf", x"f773", 
            x"ec58", x"0318", x"2499", x"28ba", 
            x"efd8", x"cac3", x"01d3", x"1b49", 
            x"e6d1", x"d8c5", x"05d0", x"032e", 
            x"d9f0", x"d727", x"eadc", x"08c5", 
            x"1dd4", x"fdc4", x"ddf5", x"f068", 
            x"15a8", x"2d31", x"279f", x"2778", 
            x"250c", x"02ac", x"f234", x"077a", 
            x"2da5", x"2a0b", x"f875", x"ec46", 
            x"029c", x"0d97", x"1e35", x"16a7", 
            x"e84e", x"ccbe", x"ea7a", x"2991", 
            x"3916", x"06d3", x"ed6f", x"051d", 
            x"0d8b", x"0972", x"0e3c", x"0eda", 
            x"eb38", x"cf0f", x"0a01", x"4b1f", 
            x"313d", x"d79a", x"cc89", x"1544", 
            x"1ffa", x"eb56", x"e4d2", x"2059", 
            x"3ba6", x"0936", x"f00e", x"1a2c", 
            x"334a", x"2381", x"1c1a", x"329e", 
            x"45af", x"2e32", x"1cc5", x"3a6e", 
            x"3f74", x"1d62", x"f932", x"df71", 
            x"efd0", x"0a42", x"0208", x"ee4f", 
            x"e8ae", x"f3a0", x"0a00", x"1e47", 
            x"0eb3", x"f4a7", x"ed1d", x"ed5c", 
            x"e749", x"d42e", x"c9fc", x"ed22", 
            x"0457", x"ef9f", x"d4f5", x"df5e", 
            x"ee52", x"def6", x"e573", x"20d6", 
            x"3add", x"ea51", x"a61a", x"e9d0", 
            x"5b46", x"463e", x"d234", x"b610", 
            x"f631", x"13ba", x"1236", x"2142", 
            x"0f26", x"d9bf", x"c07a", x"eb7c", 
            x"2536", x"0fba", x"bc66", x"995b", 
            x"d521", x"26af", x"20ff", x"e129", 
            x"e29f", x"0cc3", x"0c5e", x"d8a7", 
            x"cbf7", x"08a8", x"2b91", x"0498", 
            x"d09b", x"d496", x"ffb5", x"18a3", 
            x"00d1", x"c91d", x"c1ff", x"fe22", 
            x"144d", x"eef4", x"d3c8", x"e503", 
            x"0aef", x"01e5", x"d754", x"d82c", 
            x"df95", x"d319", x"cee9", x"c36c", 
            x"bf16", x"e509", x"1d1a", x"2e83", 
            x"030a", x"df49", x"017c", x"2153", 
            x"ec14", x"b9fc", x"e26b", x"296a", 
            x"2b78", x"ebfe", x"cbb4", x"f3e1", 
            x"1dd2", x"006b", x"dcb5", x"ea60", 
            x"0b5e", x"0ca8", x"f4e5", x"e8ea", 
            x"01a2", x"f002", x"b353", x"de9b", 
            x"2109", x"e3c1", x"8cb4", x"9d83", 
            x"e0dd", x"006d", x"f952", x"f196", 
            x"12b4", x"0cfe", x"dd28", x"efcc", 
            x"20da", x"0e0c", x"db98", x"e357", 
            x"19db", x"2a2f", x"111a", x"0488", 
            x"098b", x"3164", x"3b0b", x"0f76", 
            x"e3a0", x"dee3", x"0434", x"1582", 
            x"163b", x"18b9", x"036a", x"005d", 
            x"2cc4", x"4b64", x"48f2", x"23d7", 
            x"0cd4", x"1cbd", x"0e4b", x"f29a", 
            x"0dc3", x"1fd1", x"010f", x"e75b", 
            x"0b10", x"4aac", x"34cc", x"d0d9", 
            x"c3ce", x"055a", x"1498", x"0746", 
            x"05d8", x"f538", x"e7e0", x"e5b8", 
            x"f771", x"230b", x"3127", x"f443", 
            x"e405", x"1912", x"1cd9", x"0b2f", 
            x"0d99", x"3177", x"4476", x"0df1", 
            x"d5b9", x"e231", x"0b43", x"1df5", 
            x"25fc", x"2964", x"3230", x"1f8d", 
            x"e955", x"dfe8", x"0f7f", x"463f", 
            x"4bb0", x"01ee", x"ce84", x"fbda", 
            x"2d4e", x"21aa", x"0b25", x"e753", 
            x"c705", x"f0ff", x"2b80", x"fc0d", 
            x"adb5", x"c2c7", x"3171", x"5ab8", 
            x"1fd0", x"f832", x"0188", x"0534", 
            x"06ac", x"2448", x"21e9", x"f4fa", 
            x"d4ea", x"0887", x"4e49", x"2041", 
            x"ca19", x"ec19", x"3df2", x"225c", 
            x"c948", x"c381", x"f639", x"1181", 
            x"1980", x"0762", x"0285", x"1b45", 
            x"25f6", x"295b", x"2614", x"00a4", 
            x"f8fe", x"1c3e", x"1c85", x"047d", 
            x"f54d", x"c9ad", x"bad8", x"efce", 
            x"219b", x"144d", x"d789", x"b65f", 
            x"d210", x"0e6a", x"251f", x"11ee", 
            x"e639", x"d941", x"16df", x"4b6c", 
            x"3029", x"ff91", x"13dd", x"409a", 
            x"33ae", x"19b1", x"2322", x"16fe", 
            x"f25a", x"db8e", x"f794", x"193d", 
            x"10e4", x"fd97", x"ebc1", x"dceb", 
            x"e7c2", x"1082", x"1e4f", x"ffe1", 
            x"ef00", x"efaa", x"de8f", x"d8f5", 
            x"facb", x"0d45", x"e5e9", x"cda1", 
            x"cd18", x"ef18", x"350b", x"2a5d", 
            x"d62b", x"d953", x"0fb4", x"f3da", 
            x"e418", x"18e3", x"21d4", x"000a", 
            x"f481", x"f850", x"1645", x"30b9", 
            x"143f", x"f614", x"0821", x"1e3c", 
            x"17f6", x"2884", x"4876", x"3697", 
            x"3290", x"4018", x"20ee", x"fc32", 
            x"effc", x"f859", x"ffc1", x"f052", 
            x"f7f8", x"ee09", x"d41d", x"edb2", 
            x"1699", x"1fed", x"10ac", x"14ec", 
            x"155c", x"0bea", x"0566", x"f51a", 
            x"ea10", x"0e9c", x"1aae", x"f78b", 
            x"fa79", x"1629", x"11cd", x"103b", 
            x"2831", x"3842", x"4581", x"2417", 
            x"df7d", x"cc48", x"f6eb", x"17dd", 
            x"1c80", x"3384", x"3bd6", x"1335", 
            x"071a", x"20e4", x"21de", x"0c68", 
            x"f7db", x"e207", x"dc61", x"ed1e", 
            x"eb61", x"eb6c", x"f592", x"efe2", 
            x"0389", x"1c57", x"1679", x"f8fb", 
            x"dc02", x"dc6e", x"e60b", x"fdde", 
            x"fb7d", x"e267", x"d323", x"c932", 
            x"d8ed", x"0745", x"17b4", x"e8a6", 
            x"c1e3", x"d1a5", x"e065", x"dfd0", 
            x"e3e9", x"db9f", x"d234", x"c7c0", 
            x"bb38", x"c031", x"e680", x"fdca", 
            x"fdb7", x"0788", x"fa3c", x"ff19", 
            x"3c16", x"4845", x"fcfe", x"f00e", 
            x"23ff", x"3f26", x"33a8", x"1916", 
            x"fd35", x"f5f6", x"0d3b", x"20d5", 
            x"0d11", x"d34f", x"e9ad", x"2e45", 
            x"3545", x"16c0", x"2132", x"16e9", 
            x"e35e", x"f4ff", x"0e49", x"de68", 
            x"bf46", x"ee82", x"1b0e", x"2ed3", 
            x"0c2a", x"dd7d", x"ef78", x"1633", 
            x"282f", x"0eda", x"e7c8", x"d8dc", 
            x"f9c8", x"0bed", x"ea2f", x"e07e", 
            x"17b2", x"3b59", x"1c8a", x"e1cd", 
            x"d736", x"0086", x"176c", x"f677", 
            x"ee88", x"05b9", x"f7b3", x"d3fa", 
            x"cde7", x"d95b", x"e4f4", x"09a4", 
            x"1b42", x"f1a8", x"c601", x"c2ed", 
            x"b7e5", x"c4a0", x"ec7c", x"fab0", 
            x"e652", x"cb53", x"ab24", x"a21f", 
            x"c116", x"eaa9", x"0dc2", x"ff86", 
            x"d786", x"c79c", x"e25f", x"071b", 
            x"0f0c", x"07f0", x"f752", x"f193", 
            x"0978", x"1d6e", x"0000", x"dea2", 
            x"f3d3", x"1ab1", x"2c99", x"1cae", 
            x"0c21", x"2168", x"32f2", x"1b78", 
            x"ec66", x"d86d", x"f61b", x"fa63", 
            x"d898", x"e34c", x"0e4f", x"1efe", 
            x"2a00", x"08b0", x"d6ac", x"e084", 
            x"fd82", x"fbe8", x"1830", x"13bc", 
            x"b60e", x"82a5", x"ae09", x"df70", 
            x"e5d0", x"e2ac", x"d4fa", x"d130", 
            x"d7f9", x"eb8e", x"fefb", x"1635", 
            x"fc22", x"dad0", x"f94b", x"1033", 
            x"f677", x"f90b", x"0676", x"0417", 
            x"116f", x"160f", x"331e", x"4c2d", 
            x"1e89", x"ed81", x"155c", x"510c", 
            x"512a", x"0b56", x"d132", x"09e7", 
            x"6396", x"4b50", x"f62b", x"016e", 
            x"420b", x"2766", x"fea9", x"0241", 
            x"f2a8", x"f13c", x"f7f0", x"e3d5", 
            x"fb3c", x"136f", x"ec12", x"d154", 
            x"d27c", x"ce0b", x"c6cc", x"ca5c", 
            x"cae3", x"d1f6", x"e7cf", x"034d", 
            x"0496", x"086d", x"35b4", x"3557", 
            x"f2ba", x"c558", x"f46d", x"2e9f", 
            x"1f3c", x"0178", x"1398", x"3807", 
            x"2b96", x"1b1d", x"4e58", x"610d", 
            x"1acf", x"fcf2", x"2930", x"3b4e", 
            x"0644", x"dd25", x"1651", x"4c1e", 
            x"25b1", x"013a", x"0160", x"ebc6", 
            x"df65", x"1151", x"3943", x"1873", 
            x"fd8e", x"082f", x"f2db", x"e7ef", 
            x"fa4f", x"0fca", x"f8ed", x"da75", 
            x"f47e", x"0f1f", x"f5db", x"dc9f", 
            x"fe48", x"2524", x"2c9a", x"166d", 
            x"0222", x"d024", x"b8f0", x"055f", 
            x"5299", x"2181", x"b983", x"91eb", 
            x"c987", x"f9e7", x"f6d8", x"edfc", 
            x"e12c", x"dd16", x"f24e", x"fe0e", 
            x"e26a", x"d6b9", x"0876", x"42b4", 
            x"364d", x"220a", x"2484", x"1564", 
            x"0fe2", x"3195", x"3a0c", x"218a", 
            x"0994", x"25d4", x"5106", x"3b45", 
            x"1dce", x"2b97", x"1bc0", x"1766", 
            x"3b58", x"1404", x"cd7f", x"fc2f", 
            x"3f3f", x"4510", x"249e", x"ef85", 
            x"d4e2", x"f635", x"08eb", x"d4aa", 
            x"b2ae", x"9982", x"a35d", x"dacb", 
            x"01a9", x"df09", x"af6c", x"db2d", 
            x"2140", x"206d", x"e50c", x"b23f", 
            x"c4fd", x"14b6", x"36da", x"e375", 
            x"b581", x"0485", x"323e", x"19c9", 
            x"09d4", x"04b9", x"fe5c", x"e0e2", 
            x"d5eb", x"279e", x"4c27", x"ee5e", 
            x"d377", x"11ac", x"30c4", x"20e9", 
            x"0542", x"f5bc", x"f393", x"ef53", 
            x"ef70", x"054b", x"0892", x"e30d", 
            x"ec34", x"f8eb", x"e28e", x"eb4b", 
            x"fd36", x"e9b7", x"d7a5", x"f1bc", 
            x"1ba7", x"0229", x"d627", x"0b78", 
            x"36dd", x"f2f7", x"c562", x"f65c", 
            x"23bd", x"2320", x"efe7", x"d77f", 
            x"171e", x"475b", x"328d", x"3852", 
            x"48d9", x"2358", x"0f69", x"1ab0", 
            x"0da6", x"1991", x"4e13", x"45c0", 
            x"040c", x"f375", x"0d75", x"fa0c", 
            x"f1ba", x"0a0c", x"e21c", x"b572", 
            x"d491", x"0261", x"01ed", x"cfe5", 
            x"af1e", x"ea29", x"3000", x"15fa", 
            x"e2e4", x"f007", x"f9f7", x"eb48", 
            x"21e3", x"426c", x"3365", x"306f", 
            x"13e2", x"eef6", x"0e41", x"23aa", 
            x"e2da", x"f9fc", x"53ac", x"18a9", 
            x"bc3e", x"008a", x"4b7f", x"3184", 
            x"043f", x"ffe0", x"3161", x"4755", 
            x"15b8", x"0207", x"234c", x"18d0", 
            x"0378", x"1585", x"1694", x"f09a", 
            x"e4e0", x"f5bf", x"e39d", x"b692", 
            x"c40f", x"09c6", x"f7d9", x"b11c", 
            x"dc94", x"fd35", x"d122", x"eaae", 
            x"2a9c", x"2ab3", x"ed92", x"df83", 
            x"185e", x"337b", x"0732", x"d499", 
            x"c261", x"c5ab", x"ebc9", x"15b2", 
            x"0518", x"cec8", x"cc48", x"f74a", 
            x"023d", x"dec3", x"f800", x"263d", 
            x"00f5", x"e157", x"ffb9", x"030d", 
            x"f641", x"f90a", x"f7e3", x"fa15", 
            x"ce91", x"e130", x"302d", x"3589", 
            x"17c4", x"1407", x"e8d8", x"ccc2", 
            x"0403", x"3cae", x"292f", x"ce93", 
            x"b66e", x"e618", x"2af2", x"1df4", 
            x"eae8", x"cf55", x"b564", x"d31b", 
            x"2797", x"2f7b", x"bb3a", x"9165", 
            x"fc57", x"58ee", x"0277", x"ad42", 
            x"eb3e", x"3016", x"114e", x"dd5a"
        ),
        -- Block 1
        (
            x"f10d", x"263d", x"2d0e", x"fe9c", 
            x"f3a0", x"f5f5", x"ee8b", x"f77a", 
            x"082b", x"f4a7", x"ddd1", x"ed21", 
            x"e5c6", x"eb9b", x"e71b", x"dcdb", 
            x"fda1", x"09dc", x"03f0", x"fa72", 
            x"e92a", x"e9a1", x"1e70", x"3401", 
            x"271a", x"07f2", x"e14d", x"1309", 
            x"56ac", x"2cae", x"0d0b", x"249e", 
            x"23e0", x"422b", x"4bfc", x"06b7", 
            x"f1d9", x"2faa", x"403c", x"2c79", 
            x"ec61", x"d549", x"104a", x"1dd1", 
            x"0205", x"fdfd", x"13e7", x"0a0b", 
            x"ebb4", x"fa44", x"05d7", x"0bc3", 
            x"160c", x"f07e", x"ca0f", x"f93a", 
            x"f13a", x"bb6b", x"fa56", x"2ba6", 
            x"ef01", x"a95e", x"a769", x"d02a", 
            x"fddf", x"ea0e", x"b7e5", x"d2fd", 
            x"1f63", x"3b60", x"03bf", x"bc7e", 
            x"d0f1", x"0884", x"f80c", x"e6aa", 
            x"ead9", x"efb0", x"11d9", x"2302", 
            x"1274", x"1bfb", x"2d33", x"1aa4", 
            x"0052", x"fd14", x"05b5", x"26ec", 
            x"1296", x"d2ac", x"ea60", x"166e", 
            x"04eb", x"ee02", x"f2bd", x"e674", 
            x"e096", x"e41c", x"03c3", x"151f", 
            x"f3d4", x"e424", x"d061", x"d79e", 
            x"e931", x"d6f8", x"f36b", x"3029", 
            x"1446", x"f4bb", x"076e", x"f8e8", 
            x"fe41", x"0007", x"c38f", x"dce5", 
            x"2484", x"0428", x"b521", x"e82f", 
            x"58bf", x"4917", x"fada", x"f9ad", 
            x"0ce2", x"f656", x"e0c8", x"0b00", 
            x"1ef4", x"fc6d", x"016d", x"11c6", 
            x"f896", x"dc86", x"e525", x"f0ad", 
            x"d844", x"d136", x"109a", x"4db7", 
            x"4d40", x"12a6", x"0143", x"4b30", 
            x"5603", x"f953", x"f586", x"2dba", 
            x"4ede", x"6ce7", x"3c7f", x"fab1", 
            x"245c", x"553d", x"3494", x"00c3", 
            x"e3f9", x"0813", x"471c", x"3dab", 
            x"2356", x"1efa", x"158a", x"1983", 
            x"1760", x"f187", x"d474", x"dbac", 
            x"f7c7", x"fa2d", x"f3e6", x"1f68", 
            x"15a5", x"c24d", x"bb59", x"1103", 
            x"2cd5", x"d71e", x"923e", x"e51c", 
            x"4363", x"1ac4", x"db71", x"e5ef", 
            x"25e2", x"2938", x"e97e", x"e5f8", 
            x"186a", x"2900", x"05b8", x"ee98", 
            x"010f", x"0cfc", x"1b4a", x"14b0", 
            x"fa0d", x"fe38", x"0e2b", x"0723", 
            x"0eb8", x"216c", x"15ab", x"fbd1", 
            x"edef", x"f35d", x"0aa3", x"07fc", 
            x"ed11", x"ebd9", x"1e3c", x"41e1", 
            x"160f", x"eb6d", x"09ae", x"3224", 
            x"1eae", x"d33b", x"b316", x"e918", 
            x"187b", x"003c", x"dd4f", x"d442", 
            x"d171", x"cb2f", x"dcdc", x"e466", 
            x"e5a3", x"ee9b", x"ea45", x"efa8", 
            x"10ba", x"0e6a", x"f277", x"efae", 
            x"0340", x"1f78", x"1cc4", x"edd3", 
            x"ea49", x"09e1", x"01d9", x"ed8c", 
            x"ee06", x"ed42", x"c507", x"bc93", 
            x"ef44", x"f875", x"c5e7", x"999f", 
            x"b39d", x"0698", x"15f0", x"d869", 
            x"cea0", x"f50a", x"06c1", x"1734", 
            x"0b75", x"d449", x"e632", x"20bd", 
            x"1a7b", x"0ee7", x"f6e5", x"ff9e", 
            x"3cea", x"3738", x"f5f7", x"f86e", 
            x"0440", x"f635", x"087e", x"18cd", 
            x"0903", x"0efe", x"2d0a", x"19e0", 
            x"051f", x"0bdb", x"1616", x"063b", 
            x"e8d0", x"f9ad", x"1d10", x"0ca3", 
            x"f239", x"f753", x"f66c", x"0647", 
            x"f973", x"d912", x"db9d", x"0977", 
            x"0d52", x"e155", x"d038", x"cfab", 
            x"f0f6", x"f594", x"dded", x"d1e3", 
            x"fe05", x"19fd", x"e4d2", x"c562", 
            x"ecc1", x"0f3d", x"f362", x"b095", 
            x"cc54", x"1afc", x"eaf3", x"9f37", 
            x"b1e3", x"fc12", x"0793", x"e203", 
            x"dc8b", x"0a92", x"27cc", x"0515", 
            x"ea18", x"fd15", x"1144", x"07cc", 
            x"02e1", x"fac8", x"f4c6", x"1683", 
            x"2c4a", x"1d70", x"23e2", x"2ba2", 
            x"fddb", x"e7f2", x"0722", x"000f", 
            x"f050", x"1e19", x"4e21", x"1505", 
            x"d3ad", x"e2cb", x"0346", x"1058", 
            x"f8c9", x"d369", x"c591", x"c9af", 
            x"d5b2", x"d6f3", x"e6b7", x"1c5e", 
            x"13f5", x"e2ff", x"ed74", x"19a1", 
            x"3520", x"3d34", x"0fca", x"e716", 
            x"09fc", x"2382", x"0887", x"028f", 
            x"34e2", x"3ff9", x"30f5", x"3adf", 
            x"4275", x"2df6", x"17c8", x"1888", 
            x"1dd9", x"fda5", x"d13c", x"f065", 
            x"42d1", x"39a1", x"f063", x"f13a", 
            x"0a70", x"fbda", x"e231", x"f3af", 
            x"0750", x"fe0a", x"e95d", x"e366", 
            x"fd43", x"1c52", x"246a", x"1775", 
            x"fa00", x"0aaa", x"2143", x"2036", 
            x"1030", x"f676", x"f60b", x"135a", 
            x"293e", x"101b", x"feed", x"094e", 
            x"1ed7", x"258d", x"04fb", x"f2ee", 
            x"06d6", x"3d87", x"3507", x"ede2", 
            x"1a99", x"6f61", x"1b77", x"de43", 
            x"498f", x"502f", x"cf62", x"a472", 
            x"f294", x"419f", x"2a5a", x"bca5", 
            x"9270", x"e52e", x"37c5", x"1bf7", 
            x"dd66", x"c324", x"da26", x"01b4", 
            x"f70d", x"e2ab", x"f5f1", x"0b20", 
            x"04c8", x"fe09", x"f4e9", x"f4fa", 
            x"05fd", x"0d6c", x"f4ee", x"de66", 
            x"fb76", x"2023", x"0720", x"d8e1", 
            x"d865", x"1a63", x"491b", x"16a4", 
            x"ed70", x"06f5", x"15b1", x"0473", 
            x"2505", x"4aec", x"22ef", x"f168", 
            x"033d", x"37e3", x"479f", x"1a69", 
            x"fdf3", x"06b3", x"07ca", x"0c83", 
            x"1e16", x"0eca", x"e431", x"ed7e", 
            x"15fa", x"0d14", x"da7f", x"d4e4", 
            x"e5ed", x"0233", x"0074", x"e1bc", 
            x"df31", x"f5e2", x"1a18", x"214e", 
            x"f876", x"fc1b", x"1906", x"e5a1", 
            x"c348", x"0208", x"37f1", x"0d3b", 
            x"caea", x"cc70", x"0a03", x"3260", 
            x"110a", x"f4ea", x"0ec3", x"0c0f", 
            x"ef42", x"f4fe", x"fdd9", x"cf89", 
            x"cd69", x"0419", x"f41a", x"cf5e", 
            x"f15f", x"1126", x"f98d", x"00c5", 
            x"2294", x"0d5b", x"cf05", x"b80d", 
            x"e149", x"f669", x"e390", x"059d", 
            x"22ca", x"e0d8", x"e058", x"2f90", 
            x"2449", x"1583", x"19f6", x"e346", 
            x"ecb6", x"1f82", x"fefa", x"f94d", 
            x"1b67", x"114d", x"ee38", x"ecf1", 
            x"0ea5", x"16fb", x"1458", x"1454", 
            x"173f", x"085b", x"fb52", x"df0b", 
            x"d866", x"0cd3", x"02c5", x"ab75", 
            x"c523", x"f515", x"e9cc", x"07b8", 
            x"0d80", x"ec3d", x"f03d", x"f026", 
            x"f4fa", x"1084", x"ee4f", x"d35c", 
            x"e684", x"f636", x"0ed5", x"2348", 
            x"082f", x"1905", x"1e10", x"de5b", 
            x"d10d", x"101d", x"3b98", x"0aa7", 
            x"bc30", x"c75e", x"14d3", x"1df6", 
            x"07d8", x"f47a", x"f00e", x"106f", 
            x"2363", x"fb92", x"ecb9", x"176e", 
            x"359b", x"3339", x"0cfd", x"ea9a", 
            x"ef23", x"fbec", x"fb58", x"0066", 
            x"0a7c", x"e3f1", x"cd87", x"f566", 
            x"1cb4", x"012a", x"dd04", x"ecff", 
            x"ff72", x"fe77", x"e8f7", x"d639", 
            x"e22a", x"088e", x"1e81", x"010f", 
            x"c8e5", x"c2bb", x"fe6b", x"2e3b", 
            x"1dbc", x"fd0e", x"ec8e", x"fae1", 
            x"1c15", x"1967", x"fcb2", x"0acd", 
            x"1967", x"1a2d", x"fd1e", x"d2f1", 
            x"d9a3", x"0e06", x"3a99", x"3f4a", 
            x"15a0", x"ddbb", x"f123", x"2a94", 
            x"25e4", x"f4af", x"dda0", x"ea58", 
            x"ea87", x"e7d8", x"0916", x"0cce", 
            x"e198", x"dcc3", x"fd56", x"f8d4", 
            x"082e", x"03d1", x"b383", x"b716", 
            x"fc2a", x"0dbb", x"1d68", x"13d4", 
            x"ecf2", x"1be9", x"43ce", x"f995", 
            x"f188", x"361a", x"303b", x"0f01", 
            x"fc3e", x"0d6f", x"2a39", x"1dd6", 
            x"249f", x"4984", x"39a2", x"e59d", 
            x"c333", x"06bd", x"3850", x"08c3", 
            x"e921", x"1066", x"1a67", x"f0c5", 
            x"df18", x"eee0", x"0205", x"f747", 
            x"d970", x"bd12", x"bd0d", x"dc0b", 
            x"1ecf", x"405d", x"03a0", x"b151", 
            x"b783", x"f3f7", x"0f0d", x"0d54", 
            x"f0f3", x"db4e", x"eadf", x"f865", 
            x"e66a", x"e13f", x"eca1", x"0ac5", 
            x"14db", x"e3a9", x"db26", x"2071", 
            x"36f5", x"088f", x"f52e", x"e78d", 
            x"ef41", x"0782", x"0785", x"ff0d", 
            x"f2c8", x"ec26", x"fff9", x"1d57", 
            x"240b", x"11d4", x"03f3", x"0db1", 
            x"0fc1", x"070d", x"fb77", x"f76b", 
            x"edea", x"ef11", x"f3f7", x"f5a8", 
            x"fbb3", x"eb6a", x"df1d", x"fa14", 
            x"0a6e", x"f4b6", x"eae6", x"eb98", 
            x"de7b", x"d170", x"d764", x"f5c0", 
            x"0d48", x"0312", x"e30e", x"cff6", 
            x"d8f8", x"efc4", x"0168", x"1216", 
            x"17e8", x"06d3", x"ed0f", x"ff49", 
            x"2ea1", x"285d", x"ed22", x"d98b", 
            x"f533", x"1404", x"1eee", x"0504", 
            x"f59d", x"188b", x"2176", x"1cfe", 
            x"1116", x"00c7", x"05c7", x"1a5e", 
            x"1662", x"062f", x"1461", x"179b", 
            x"fe89", x"fde8", x"22a3", x"2961", 
            x"f8e5", x"d6fd", x"f8c2", x"1ae8", 
            x"1ce0", x"0711", x"f002", x"f70d", 
            x"12dc", x"166c", x"1003", x"0bce", 
            x"01df", x"ff24", x"0b9b", x"14de", 
            x"102d", x"0528", x"f9dc", x"f0bb", 
            x"1996", x"33ac", x"f440", x"c3ce", 
            x"f7d0", x"35b3", x"1722", x"e2a0", 
            x"ee30", x"1684", x"25ed", x"12c3", 
            x"07da", x"1b10", x"1e60", x"2014", 
            x"247f", x"1c7e", x"1e64", x"2ced", 
            x"1d42", x"08d0", x"164c", x"2d52", 
            x"15de", x"00ab", x"168d", x"182e", 
            x"fa43", x"ed8e", x"ffeb", x"2bdc", 
            x"2d08", x"02bc", x"fd95", x"060f", 
            x"f486", x"f6e8", x"04a1", x"eae6", 
            x"ecd2", x"037b", x"ff36", x"fea1", 
            x"0a6f", x"1c06", x"0acf", x"eab2", 
            x"f58a", x"0a7b", x"00c1", x"f33b", 
            x"f7d1", x"14ee", x"19dc", x"f708", 
            x"f6d9", x"fce8", x"1246", x"28f2", 
            x"09d3", x"eb64", x"00a7", x"19f5", 
            x"1404", x"f71d", x"ec71", x"022e", 
            x"029e", x"f59d", x"e138", x"caf0", 
            x"c672", x"e3a8", x"ff71", x"0be6", 
            x"ea9e", x"d1b2", x"e54b", x"f943", 
            x"0c5b", x"2199", x"0864", x"e0cc", 
            x"e22c", x"04ca", x"277f", x"2560", 
            x"0b2e", x"0178", x"0149", x"ffe4", 
            x"1618", x"19fd", x"ec9f", x"db21", 
            x"16f5", x"2d53", x"f904", x"db01", 
            x"f1a4", x"0abe", x"0f89", x"04c9", 
            x"faf1", x"fe74", x"095d", x"073c", 
            x"09fb", x"0f60", x"fab0", x"dceb", 
            x"d128", x"e4cd", x"f629", x"dda4", 
            x"bedd", x"d076", x"efd3", x"f02e", 
            x"d6c1", x"cc8d", x"da6e", x"f122", 
            x"e615", x"dd1b", x"0630", x"1ae0", 
            x"eb98", x"ccf6", x"ef4e", x"06ff", 
            x"dd4e", x"bdb3", x"eff3", x"0016", 
            x"e13e", x"e073", x"f269", x"01d7", 
            x"f66d", x"ef7f", x"f6bf", x"0462", 
            x"02dc", x"e936", x"f406", x"0b2c", 
            x"0434", x"f2bb", x"0578", x"0630", 
            x"d810", x"d1f3", x"eb0f", x"e067", 
            x"e5f1", x"e2d5", x"ce55", x"d353", 
            x"d6b5", x"dca5", x"e833", x"f232", 
            x"f0e1", x"e30f", x"d270", x"ddd2", 
            x"f2d2", x"f657", x"e65a", x"e4c5", 
            x"041b", x"1003", x"05be", x"fee4", 
            x"fc97", x"1cdd", x"2f8b", x"feb2", 
            x"ea55", x"0dad", x"28cb", x"1269", 
            x"edc3", x"ee5c", x"0147", x"f950", 
            x"06b3", x"1519", x"f5d9", x"d03e", 
            x"e69c", x"1653", x"1c23", x"fce3", 
            x"e625", x"f862", x"179a", x"203d", 
            x"f99c", x"f053", x"f86e", x"f8e5", 
            x"179b", x"357b", x"097c", x"e104", 
            x"0b02", x"3925", x"3a1a", x"1f00", 
            x"f60d", x"07c5", x"4ef1", x"49c2", 
            x"10ea", x"0aaf", x"2986", x"3c25", 
            x"3b7c", x"2286", x"10f9", x"0ffd"
        ),
        -- Block 0
        (
            x"095e", x"0b10", x"1c72", x"176f", 
            x"ffc4", x"ea06", x"0d3f", x"2699", 
            x"072b", x"f936", x"00d1", x"0f2b", 
            x"0e6d", x"e9ef", x"d74f", x"02b5", 
            x"1b5a", x"f931", x"dae5", x"f192", 
            x"16f5", x"3915", x"3d10", x"2220", 
            x"f5bd", x"fc22", x"3f54", x"5108", 
            x"3804", x"2aae", x"20e1", x"134e", 
            x"3188", x"5c82", x"4dc3", x"02ad", 
            x"d9db", x"021b", x"2ae3", x"3e8e", 
            x"1cc8", x"e820", x"d691", x"e390", 
            x"0a7c", x"1803", x"f306", x"e961", 
            x"e983", x"d8ae", x"d06a", x"dcba", 
            x"fdd7", x"03c1", x"f35f", x"d540", 
            x"c0ad", x"daf0", x"f82d", x"02af", 
            x"fe62", x"f07c", x"eee2", x"ed95", 
            x"f346", x"13f5", x"21c7", x"076d", 
            x"fcd0", x"1291", x"1f0f", x"f724", 
            x"ec55", x"1f9a", x"29e9", x"054e", 
            x"05fc", x"2ab4", x"2767", x"037a", 
            x"166a", x"4cca", x"3330", x"f142", 
            x"0048", x"1b1d", x"0b61", x"fe47", 
            x"02e2", x"04d7", x"f633", x"ea33", 
            x"f469", x"f2bd", x"dff8", x"ed48", 
            x"fcc5", x"f9df", x"eb35", x"df7a", 
            x"f683", x"0641", x"e657", x"df5b", 
            x"f3fe", x"f6cb", x"ecc5", x"dcaa", 
            x"f04d", x"10d3", x"fde3", x"f010", 
            x"081f", x"08d0", x"dfc0", x"e357", 
            x"10a5", x"15e5", x"e33a", x"bf2c", 
            x"f745", x"26a3", x"03b9", x"e447", 
            x"fd75", x"0853", x"eaa7", x"e45b", 
            x"fd69", x"feb3", x"f732", x"06b8", 
            x"eb45", x"b826", x"d0f1", x"03f6", 
            x"f7fa", x"d65b", x"d850", x"f8b7", 
            x"f424", x"ef45", x"16a0", x"25df", 
            x"115b", x"e79e", x"e7b6", x"1889", 
            x"1973", x"0264", x"1272", x"0932", 
            x"f58b", x"191e", x"3c26", x"3d81", 
            x"26e9", x"fddf", x"fe51", x"28f3", 
            x"2815", x"0145", x"e8ba", x"0d64", 
            x"3740", x"2ca4", x"008b", x"e2a9", 
            x"f2d3", x"2205", x"1b5a", x"e7d3", 
            x"d47a", x"d5b1", x"dbe9", x"f14d", 
            x"fffb", x"e3dc", x"ccae", x"f335", 
            x"0375", x"df33", x"e57b", x"f321", 
            x"d67d", x"cf50", x"efbc", x"02a4", 
            x"05d6", x"040a", x"fc69", x"16d8", 
            x"1d21", x"fc6f", x"fc9c", x"0cbf", 
            x"ec30", x"e50d", x"1a7a", x"13dc", 
            x"de39", x"e712", x"1713", x"0d61", 
            x"f00d", x"f7bc", x"f6ce", x"dfa5", 
            x"e276", x"f928", x"f307", x"ecc8", 
            x"f7e3", x"0958", x"098b", x"f1ff", 
            x"e2a2", x"fe9c", x"1331", x"1365", 
            x"0a18", x"f4f2", x"f78a", x"0a72", 
            x"182c", x"1c37", x"1273", x"18dc", 
            x"201f", x"fea3", x"f2fb", x"1e0e", 
            x"35e8", x"0fb2", x"f39b", x"117a", 
            x"3202", x"3058", x"166f", x"fcb5", 
            x"fd4a", x"182f", x"31bb", x"27c6", 
            x"f6ff", x"d76d", x"f25e", x"1376", 
            x"03a5", x"e1e4", x"e7be", x"fd97", 
            x"ff7c", x"04e5", x"0f88", x"02dc", 
            x"f3dc", x"f903", x"0903", x"0530", 
            x"e395", x"dedf", x"f74e", x"f26b", 
            x"e5d3", x"e622", x"f17a", x"11cc", 
            x"0313", x"e0f5", x"f7b5", x"1403", 
            x"f5b7", x"e14a", x"fe16", x"1e7c", 
            x"1bb8", x"0f59", x"06cd", x"f90e", 
            x"ffae", x"122e", x"17e0", x"0938", 
            x"1252", x"235c", x"1fb6", x"0061", 
            x"e9a4", x"09fa", x"219a", x"04b0", 
            x"f7bb", x"f6ac", x"f92b", x"0b20", 
            x"13d1", x"041c", x"f1d3", x"e909", 
            x"f03f", x"08c1", x"fbf0", x"e44d", 
            x"e097", x"df2c", x"ed86", x"0006", 
            x"f127", x"cb53", x"b229", x"c834", 
            x"f839", x"094f", x"e936", x"f3c5", 
            x"06c5", x"d50e", x"ac60", x"e311", 
            x"3d67", x"1be2", x"c056", x"a3ca", 
            x"d09f", x"11b7", x"2c5b", x"f4a7", 
            x"d9d2", x"06a5", x"09b8", x"f4ee", 
            x"fbcc", x"050b", x"e8ff", x"f413", 
            x"253b", x"0d10", x"d9dc", x"eb91", 
            x"f993", x"f749", x"0592", x"091c", 
            x"0821", x"f0a1", x"d10f", x"d6b6", 
            x"0660", x"37e5", x"28fc", x"e0d6", 
            x"ddc6", x"2367", x"323b", x"0456", 
            x"045d", x"2ddd", x"362d", x"1000", 
            x"067e", x"2e35", x"4a25", x"29e7", 
            x"18d9", x"3518", x"09d2", x"dbc4", 
            x"0890", x"438b", x"48df", x"1370", 
            x"04f9", x"2270", x"0939", x"ea57", 
            x"df7f", x"dae2", x"eb7e", x"0713", 
            x"0c37", x"ed13", x"cad5", x"d083", 
            x"0a18", x"34c0", x"1ef7", x"c414", 
            x"8fdb", x"c962", x"06d7", x"ee42", 
            x"c04c", x"ca8c", x"fb6e", x"1171", 
            x"f621", x"e19a", x"df01", x"d8d1", 
            x"f318", x"4e21", x"64d9", x"f6f1", 
            x"b292", x"f2ba", x"4265", x"2d34", 
            x"ed5c", x"f47b", x"1426", x"0add", 
            x"1646", x"157c", x"f749", x"fc2e", 
            x"ffdc", x"0a8f", x"1333", x"073f", 
            x"f6ef", x"e0cf", x"d0e4", x"0cfa", 
            x"24f3", x"e778", x"d049", x"f78f", 
            x"1785", x"065f", x"ebef", x"1407", 
            x"2dd0", x"efa9", x"f191", x"2877", 
            x"25a6", x"1adb", x"1fc9", x"27ff", 
            x"0cb6", x"fadb", x"04d0", x"1c31", 
            x"1fa8", x"1c39", x"2291", x"0f35", 
            x"f80d", x"ddb0", x"13eb", x"70b8", 
            x"3675", x"dc1c", x"e895", x"243e", 
            x"4bdc", x"3b00", x"245d", x"052a", 
            x"0e87", x"3935", x"4c67", x"16ab", 
            x"0394", x"23e7", x"3683", x"3975", 
            x"1a60", x"0b9b", x"2593", x"1bb1", 
            x"fdc7", x"01a4", x"f114", x"fbed", 
            x"12ea", x"14f4", x"e0f1", x"c802", 
            x"f0bf", x"f756", x"f366", x"fda3", 
            x"e8e9", x"c687", x"dcef", x"dfc5", 
            x"e219", x"f651", x"041f", x"f14c", 
            x"dcbc", x"ebb1", x"ff2b", x"fe00", 
            x"f414", x"ee78", x"e84a", x"f380", 
            x"ff0f", x"0d6b", x"14d6", x"f1d7", 
            x"e694", x"fa56", x"fe4c", x"fe48", 
            x"1241", x"2ae4", x"159f", x"e9aa", 
            x"e38c", x"0bed", x"246c", x"2100", 
            x"14af", x"079b", x"e720", x"de0f", 
            x"f5c1", x"0cc0", x"0ac9", x"f867", 
            x"f4b7", x"f811", x"f14a", x"fc45", 
            x"14aa", x"097b", x"f03a", x"eedb", 
            x"ef35", x"f2d6", x"007a", x"f606", 
            x"dc39", x"d29f", x"e697", x"0556", 
            x"03f3", x"e16f", x"c9e3", x"d49c", 
            x"f7a8", x"07a4", x"ef70", x"dab2", 
            x"ea5f", x"f400", x"e883", x"eaba", 
            x"ff0d", x"0904", x"fd35", x"e82b", 
            x"ebd7", x"fe95", x"fcae", x"04b7", 
            x"0bb3", x"ff40", x"00f8", x"0dff", 
            x"06e7", x"f24a", x"fad5", x"08f1", 
            x"0543", x"f747", x"fa4b", x"1bc4", 
            x"22fe", x"0cc6", x"112d", x"1eb0", 
            x"0c19", x"fbea", x"12c1", x"1c09", 
            x"022f", x"f7e6", x"f98d", x"f6c0", 
            x"ed9d", x"f370", x"0a3d", x"fd5d", 
            x"d6aa", x"d810", x"f51a", x"f7df", 
            x"ef9f", x"e67d", x"e0e8", x"ee4b", 
            x"f7b0", x"eb1d", x"de83", x"e8a0", 
            x"eed0", x"f3ee", x"f8fa", x"f4f0", 
            x"fadf", x"fffd", x"ede4", x"f458", 
            x"0910", x"fff7", x"ec76", x"f58f", 
            x"0c52", x"172b", x"1b25", x"05e3", 
            x"ef69", x"00ca", x"1b7e", x"1a94", 
            x"0dfb", x"fa39", x"efb7", x"f97b", 
            x"11d3", x"2795", x"1729", x"f510", 
            x"0006", x"17e4", x"10e8", x"fd5e", 
            x"05cb", x"16d1", x"03a9", x"f453", 
            x"04c2", x"05a8", x"f30a", x"ed31", 
            x"01f8", x"0ee2", x"f362", x"eb8b", 
            x"065f", x"0caf", x"f862", x"f08b", 
            x"02b9", x"08d0", x"07aa", x"19d5", 
            x"1abf", x"fe67", x"f645", x"ff17", 
            x"02bb", x"0470", x"026c", x"f12e", 
            x"eeb0", x"f581", x"ea39", x"ea8f", 
            x"f9dd", x"1019", x"1dab", x"f0f7", 
            x"c1f9", x"d5ec", x"f339", x"fc64", 
            x"0630", x"1c35", x"101d", x"d78f", 
            x"df2e", x"19c0", x"2604", x"0031", 
            x"eba7", x"f457", x"005a", x"f7b8", 
            x"fa90", x"13dc", x"0bde", x"d95a", 
            x"ddec", x"15e3", x"2a9c", x"0fb9", 
            x"fa4e", x"0323", x"09fa", x"136f", 
            x"2130", x"1346", x"fe24", x"17fc", 
            x"2a4d", x"1cd8", x"0e6a", x"0e8c", 
            x"1624", x"1f93", x"1576", x"07b3", 
            x"00e5", x"f668", x"ff27", x"0f59", 
            x"0baa", x"03c7", x"0756", x"f782", 
            x"fbce", x"12d6", x"1314", x"f369", 
            x"eb86", x"0440", x"177f", x"137a", 
            x"08b9", x"052a", x"0553", x"ef1b", 
            x"ec70", x"0737", x"048a", x"e599", 
            x"f68e", x"06fe", x"f67c", x"f4a8", 
            x"f6a1", x"05ac", x"2d34", x"126d", 
            x"df14", x"f327", x"1168", x"0dba", 
            x"0281", x"1280", x"0a73", x"e2e0", 
            x"e9f0", x"054a", x"04da", x"0de8", 
            x"0afc", x"ef91", x"ed83", x"0645", 
            x"141e", x"0bd4", x"f6ba", x"f53d", 
            x"fd92", x"eef4", x"fa6f", x"1159", 
            x"128a", x"fe7c", x"ed08", x"ee18", 
            x"f398", x"032f", x"0f65", x"08a6", 
            x"ffa9", x"f4a2", x"f4ba", x"068d", 
            x"1117", x"0203", x"006d", x"0202", 
            x"fc38", x"0380", x"03e3", x"0391", 
            x"01ba", x"06cd", x"00a3", x"ec30", 
            x"eaea", x"f686", x"f2b4", x"eada", 
            x"f4ca", x"fa8b", x"f99b", x"f445", 
            x"f01a", x"f01f", x"f3f6", x"e980", 
            x"e9d9", x"febc", x"0072", x"e59f", 
            x"dc4e", x"eeb0", x"f6a9", x"00da", 
            x"0ce8", x"f7e0", x"d6b7", x"d614", 
            x"ee1a", x"065e", x"fe12", x"ee58", 
            x"f3c7", x"edeb", x"ef0e", x"0590", 
            x"0169", x"04a9", x"0a2a", x"0105", 
            x"f0df", x"edc4", x"fa2a", x"06e3", 
            x"0df5", x"03c1", x"0420", x"0c91", 
            x"f779", x"eceb", x"0dec", x"1bfe", 
            x"07b6", x"f915", x"f9be", x"01b3", 
            x"00f9", x"020d", x"07ba", x"f7c2", 
            x"f01b", x"01af", x"065b", x"0107", 
            x"ff35", x"f953", x"f4c7", x"fb47", 
            x"0f0f", x"1417", x"fa20", x"f29a", 
            x"fe6a", x"0189", x"0300", x"0353", 
            x"faba", x"026c", x"0aec", x"fe09", 
            x"ff7b", x"0d1e", x"03a8", x"f445", 
            x"f3e6", x"038e", x"0e88", x"0186", 
            x"f624", x"f85a", x"0fed", x"15f1", 
            x"f6d6", x"fcd3", x"0e05", x"f9e7", 
            x"fc02", x"0c59", x"06c9", x"f612", 
            x"fd48", x"fca7", x"f2d9", x"fb8c", 
            x"ffae", x"011d", x"0115", x"fe77", 
            x"0f9a", x"22f8", x"144d", x"fcef", 
            x"033f", x"1e85", x"0d52", x"ee0b", 
            x"0383", x"0f47", x"13fb", x"1bc7", 
            x"028c", x"f6c7", x"15a3", x"308f", 
            x"2c3a", x"11e2", x"0205", x"08ec", 
            x"08ba", x"0707", x"08f1", x"0c69", 
            x"00a7", x"0a58", x"156d", x"030e", 
            x"fa7e", x"1595", x"1489", x"ff4f", 
            x"0105", x"056a", x"0126", x"13f5", 
            x"0ed9", x"ed35", x"0046", x"04e7", 
            x"f38d", x"e200", x"ed22", x"efef", 
            x"f67a", x"0293", x"fc74", x"e624", 
            x"f6f0", x"061b", x"00e1", x"f8c9", 
            x"0806", x"ff9f", x"f8b5", x"0914", 
            x"f618", x"eb9f", x"08b9", x"f57f", 
            x"e47b", x"fe3d", x"feb2", x"0435", 
            x"fbde", x"fa3e", x"ea0f", x"0430", 
            x"0d31", x"021c", x"038a", x"13e4", 
            x"06af", x"fc79", x"1c8b", x"2a0b", 
            x"19c6", x"0673", x"0a9e", x"0a60", 
            x"fbdd", x"19ed", x"25de", x"2205", 
            x"1797", x"0135", x"f48f", x"192e", 
            x"195f", x"fb5c", x"fada", x"f80e", 
            x"f352", x"0079", x"1206", x"fa72", 
            x"022b", x"06f0", x"fc7a", x"e89e", 
            x"f44f", x"0753", x"f817", x"ffa7", 
            x"f498", x"ea07", x"e714", x"f8d8", 
            x"0cc3", x"ffdd", x"f86a", x"f421", 
            x"eab1", x"e78b", x"effa", x"f41c", 
            x"eedd", x"ede8", x"f647", x"fef2", 
            x"fbe3", x"f46d", x"f314", x"f4a6", 
            x"f738", x"f849", x"f917", x"faa7", 
            x"fd10", x"ff04", x"0000", x"0000"
        )
    );

    -- FIFO control pointers
    signal read_p_reg, read_p_next : NATURAL;                   -- Read pointer
    
    -- Done tick
    signal done_tick_reg, done_tick_next : STD_LOGIC;
    
    -- FSM states
    type state_type is (idle, output);
    signal state_reg, state_next : state_type;
begin
    process(sysclk)
    begin
        if rising_edge(sysclk) then
            for i in 0 to n_rams-1 loop
                dout(((ir_d_width-1)+(ir_d_width*i)) downto (ir_d_width*i)) <= coeff_s(i)(read_p_reg);
            end loop;
        end if;        
    end process;
    
    -- FSM
    -- Status register
    FSM_Status : process(sysclk)
    begin
        if rising_edge(sysclk) then
            if(reset = '1') then
                state_reg <= idle;
                read_p_reg <= 0;
                done_tick_reg <= '0';
            else
                state_reg <= state_next;
                read_p_reg <= read_p_next;
                done_tick_reg <= done_tick_next;
            end if;
        end if;
    end process;
    
    -- Next state logic
    FSM_Next_state : process(state_reg, read_p_reg, start_tick)
    begin
        state_next <= state_reg;
        case state_reg is
            when idle =>
                if (start_tick = '1') then
                    state_next <= output;
                end if;
            when output =>
                if (read_p_reg = 2**bits-1) then
                    state_next <= idle;   
                end if;    
        end case;
    end process;
    
    -- Output logic
    FSM_output : process(state_reg, read_p_reg, start_tick, done_tick_reg)
    begin
        read_p_next <= read_p_reg;
        done_tick_next <= done_tick_reg;
        case state_reg is
            when idle =>
                done_tick_next <= '0';
                if (start_tick = '1') then
                    read_p_next <= 0;
                end if;
            when output =>
                if (read_p_reg = 2**bits-1) then
                    done_tick_next <= '1';
                else
                    read_p_next <= read_p_reg + 1;       
                end if;    
        end case;
    end process;
    
    -- Done tick
    done_tick <= done_tick_reg;
end Behavioral;
